-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�l�d�d�a��}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e�4�%�4��g�>���-����t/��a+��:���f�u�:�;�8�m�L���YӇ��P�'��&������_�w�}�(߁�����e9��h��U���������}���Y����^��aN�<����
�����#���Q����\��XN�N���u�%�d�8�/���������z(��c*��:���n�u�u�%�e�����Y�ƅ�5��h"��<������}�f�9� ���Y����F�G1��%���:�
�%�#�3�g�>���-����t/��=N��U���
�
�<�<�0�8�G��6����g"��x)��*�����}�d�3�*����P���F��1��!���;�
�
�
�'�+���6����g"��x)��N���u�%�a� ��0����&����|3��d:��9�������w�n�W������]ǻN��*ފ�
�<�<�2�2�l��������|3��d:��9����_�u�u������/����}F��s1��2������u�d�}�������9F���*���4��4�
�;�}�W���*����|!��d��Uʥ�c���8�9��(���Y����`2��{!��6�����u�f�w�2����I��ƹF��hX��*���<�2�0�e�6�����Y����`2��{!��6�ߊu�u�
�
��4�������)��=��*����
����u�FϺ�����O��N�������8�;���(������)��=��*����n�u�u�'�e� �������V9��N��!ʆ�������8���J�ƨ�D��^����u�
�
�
�>�4����I����E
��N��!ʆ�����]�}�W���&����^��h��U��� �u��
���(���-��� W��X����n�u�u�%�o�
��������9��h��U��� �u��
���L���YӖ��9��T��U��� �u��
���(���-���F��@ ��U���_�u�u�
�b�����&����_�!��U���
���u�l�8��Զs����Z��C��U���4�u�3�8�n�l�F���&�ƥ�l�N����� �0�����2���0����} ��N��'���n�u�u�4�#�4����:����t#��e/��:�����:�u�2�<�W�������V��E�����u�w�����������C9��Z��Y���������J���U����z(��c1��:���e�����	�1���=����5��y>��*����-�b�e�g�1�C��H߮��l/��b:��9���h�`�e�e�g�q�;���7����r4��
�����������<��W����V��{=��,����h�g����9���-Έ��VJ��d1��;����e�����3���O߮��l5��h(��M�������	�D����ƹF��X �����4�
�:�&��2����Y�Ɵ�w9��p'��O���d�n�u�u�4�3����Y����\��h�����u�u��
���W��^����F�T�����u�%��
�#�����Y�Ɵ�w9��p'��#����u�f�1� �)�W���C���V��d��Uʶ�;�!�;�u�'��(���&����F��d:��9�������w�n��������\�^�E��u�u�6�;�#�3�W���*���� 9��Z1�Oʆ�������8���Jӂ��]��G��H���d�e�n�u�w�>�����ƭ�l5��D�����f�o�����4���:����U��X����u�h�w�e�g�f�W�������R��V�����
�#�g�e�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�g�m�L���YӅ��@��CN��*���&�
�#�
�w�}�#���6����e#��x<��Eʱ�"�!�u�|�m�}�F��Y����\��V �����:�&�
�#�e�l�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��B�����D��ʴ�
�:�&�
�!�o�E��*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��X �����4�
�:�&��+�(���Y����)��t1��6���u�e�1�"�#�}�^��Y���9F������!�4�
�:�$�����J����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����4�!�4�
�8�.�(���&����`2��{!��6�����u�d�3�*����P���V��d��Uʶ�;�!�;�u�'�>�����ԓ�\��c*��:���
�����}�������	[�_�����u�:�&�4�#�<�(���
����9��N��1��������}�FϺ�����O�
N��D��u�u�6�;�#�3�W�������l
��1��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�D��w�_�u�u�8�.��������]��[�*ۖ�o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��d�e�n�u�w�>�����ƭ�l��D�����f�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��d�d�d�w�]�}�W���
������T�����f�
��o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�d�e�f�f�W�������R��V�����
�#�b�e�m��3���>����v%��eN��Cʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�w�]�}�W���
������T�����f�
��o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�d�d�g�f�W�������R��V�����
�#�
�u�w�	�(���0����p2��F����!�u�|�o�w�l�F���s���P	��C��U���6�;�!�9�c�m�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���I���9F������!�4�
�:�$�����H����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����u ��q(��U���
���
��	�%���Hӂ��]��G��H���d�d�d�d�f�l�F��H����W��_�D���_�u�u�&�0�<�W���:����^F��d:��9�������w�n��������\�^�D��u�u�4�!�>�(�ϸ�����\��PN����;�n�u�u�6�)����Ӏ��l��X
��ʺ�u�%��
�$�}�W�������@F��X ��N���u�&�2�4�w�-��������`2��C_�����u�u��
���L���Yӕ��]��V�����1�
�e�o���2���s���@��V��*ڊ�9�=�
�
�9�.���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���=�
�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��E���%�4��4��1�(���
���5��h"��<��u�u�&�2�6�}�(߁�����e9��h��*���2�o�����4��Y���9F������%�d�8�-��4�(���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����8�-��%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���@��V��*ۊ�4�
�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�F�������C9��S1�����u��
���}�J���^���F��P ��U���
�0�<�1�>�����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��G���'�:�
�'�0�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����Z��[N��G���'�:�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�E�������R��[
�����o������M���I��ƹF��^	��ʥ�`�7�!�
��3����Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*ߊ�0�4��%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���@��V��*ߊ�0�4��4��1�(���
���5��h"��<��u�u�&�2�6�}�(ځ�����l��A�����u�u��
���W��^����F�D�����%�&�2�7�3�d�W���6����}]ǻN�����9�3�%�;�3�����*����C��R��-���
�0�
�`�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����R��^	������
�!�
�$��W���-����t/��=N��U���;�9�4�
�>�����H����q)��r/�����u�<�;�9�0�-�����ד�F9��1��*���0�o�����4�ԜY�ƿ�T����*���0�!�'�
����������c9��E��C��o������!���6���F��@ ��U���_�u�u�<�9�1��������G��h=��4���4�0�4�������O����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʠ�
�:�0�!�%��!���	����G��g1�����c�b�o����0���/����aF�
�����e�n�u�u�$�:����)¹��U��W��D��������4���Y����W	��C��\�ߊu�u�<�;�;��F�������T�=��*����
����u�DϺ�����O��N�����4�u��9��2�(���	����U��V��G��������4���Y����\��XN�N���u�&�2�4�w���������\��1����e�o�����4���:����W��X����n�u�u�&�0�<�W���
����@��d:��ي�&�
�u�u���8���B�����Y�����<�
�1�
�d�}�W���5����9F������&�9�!�%�>�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʦ�9�!�%�<�%�:�A��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����;�
�
� �d�o����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���g�<�3�
�e��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����
�
�0�
�n�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������Y��*���
�e�u�u���8���&����|4�N�����u�|�_�u�w�4����	����9��h��*��u�u��
���(���-��� W��X����n�u�u�&�0�<�W�������lQ��T��!�����
����_�������V�=N��U���;�9�!�%�a�����K����`2��{!��6�����u�e�3�*����P���F��P ��U���
�
�
� �d�k����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���
�0�
�g�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������R��1�����0�
� �a�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��V ��D���9�:�0�
�2��D���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��<�����4�9�/�'�$�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʇ�;�0�
�9��8��������F��d:��9�������w�m��������l�N�����u�'�
�!��/�;���&�ߓ�l��h_�� ���m�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Z��D��&���!�
�&�
�w�}�#���6����9F������4�
�<�
�3��A���Y����v'��=N��U���;�9�4�'�;���������
9��R1��F���
�m�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��C1�����:�
�l�g�2�m�B���&����CU�=��*����
����u�FϺ�����O��N�����4�u�'�
�#���������lT��h_��*���`�c�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƭ�A9��h(��*���%�d�
�
���(���O�֓� F��d:��9�������w�n�W������]ǻN�����9�4�'�9��2�(���	����9��1�����g�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӂ��l ��h��*���g�l�4�
�#�/�W���-����t/��=N��U���;�9�2�%�1�m��������
9��h���������W�W���������h��*���
� �g�l�6�����Y�Ɵ�w9��p'�����u�<�;�9�0�-�����ד�F9��1��*���=�
�
�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��1��D���
�c�
�;�:�%�E���Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
�
�
�
�"�o�N���&����lV��T��!�����
����_������\F��d��Uʦ�2�4�u�'���(���&����_��G1�����
�u�u����>���<����N��
�����e�n�u�u�$�:��������9��1��*��
�%�'�!�%��W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����3�d�3�
�a���������F��d:��9�������w�n�W������]ǻN�����9�2�%�3�g�;�F���&����R��R����o������!���6�����Y��E��u�u�&�2�6�}����&ù��9��h\�*���6�u�u����>��Y����Z��[N��*������0�:�i�(���&����Q��N��1��������}�D�������V�=N��U���;�9�6�
���6�������9��1����g�o�����4���:����U��S�����|�_�u�u�>�3�Ͽ�����u	��{��*���g�0�e�c�%�:�E��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����!��'��8��N����ד�V��V��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�;��3���+����^9��h��*���
�f�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����}"��v<�����a�
�
�
�2��C���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*����'��:������L����`2��{!��6�����u�d�3�*����P���F��P ��U���
�
�
�
��(�E�������R��V�����
�0�u�u���8���Y���A��N�����4�u�
�
�"�o�N���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����3�
�b�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W�������	��a1�����&�<�;�3��o�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����!��'��8��A�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�
��(�E���	����`2��{!��6�����u�c�w�2����I��ƹF��^	��ʡ�%�3�
�b��l�Mύ�=����z%��r-��'���c�1�"�!�w�t�}���Y����R
��Z��A���
�m�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƾ�U�� Z��G��������4���Y����\��XN�N���u�&�2�4�w���������Z9��hZ�*��o������!���6�����Y��E��u�u�&�2�6�}����
����9��hZ�*��o������!���6�����Y��E��u�u�&�2�6�}����J����F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�����L¹��lR��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�#�-�Aځ�����l��N��1��������}�GϺ�����O��N�����4�u�8�
�c�4����Mƹ��\��c*��:���
�����}�������9F������6�'�,�3��h�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��FҊ�
�
� �a�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��@���3�
�c�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����W��C�����&�3�
�`��n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��P �����!�<�3�
�o��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��G1�*���:�2�;�<�>�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʻ�2�&�6�;�#�4����A˹��\��c*��:���
�����}�������9F������%�f�
�0�8�:��������l ��^�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�?��������l��h�� ��a�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������A��B1�F���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l ��^�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�-�!���&����^��^1��*��
�f�o����0���/����aF�N�����u�|�_�u�w�4����	����9��Q��Gڊ�f�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�/����@9��h[�*��o������!���6���F��@ ��U���_�u�u�<�9�1����*����F��B�����f�
� �`�a�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�f��(���&����W��N�&���������W��Y����G	�UךU���<�;�9�4�%�1�(���&����lW��1��E���3�
�`�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��3����:�
�l�e�8�G���&����CU�=��*����
����u�FϺ�����O��N�����4�u�'�
�#���������lT��h^��*���`�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƭ�A9��h(��*���%�d�
�
�����L����	F��s1��2������u�d�}�������9F������4�'�9�
�8�����Hʹ��V9��1��*��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������G9��E1�����l�g�0�d�c�;�(��&���5��h"��<������}�f�9� ���Y����F�D�����%��
�&�w�}�#���6����e#��x<��Fʱ�"�!�u�|�]�}�W�������C9��P1����b�o�����}���Y����R
��G1�����1�f�u�u���6��Y����Z��[N��*���
�1�
�b�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��j�MϜ�6����l�N�����u�%�&�2�5�9�B���Y����v'��=N��U���;�9�4�
�>�����@����|)��v ����u�:�%�;�9�}�3֚�8¢��lV��h_��&���u�%�'�u�]�}�W���Y����_�'��&������_�w�}�W���	����\��yN��1�����_�u�w�}�W���
����\��yN��1�����_�u�w�}�W�������	F��cN��1�����_�u�w�}�W�������	F��cN��1�����_�u�w�}�W�������\��b:��!�����n�u�w�}�WϷ�&����R9��aN�<����
�����#���Q����\��XN�N���u�u�u�<��<�(݁�Y�ƅ�5��h"��<������}�f�9� ���Y����F�N�����0�4�e��m��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����C9��C��*���u� �u����>���<����N��
�����e�n�u�u�w�}��������lW�!��U���
���
��	�%���Hӂ��]��G�U���u�u�4�
�2�(���Cө��5��h"��<������}�f�9� ���Y����F�N�����0� �;�f�m��#ύ�=����z%��r-��'���u�:�;�:�g�f�W���Y����C9��T��;ʆ�����~�W�W����Ư�^��R ���ߠ7�2�;�u�w�:����I����l ��X�Oʶ�8�:�0�!�:�d�F���M����U9��N�����u�4�u�_�w�}�W���	����[�V�����u�u�u�u�6�����GӇ��A��=N��U���u�%�&�4�#�`�W���&����U9��Q��Cӊ�%�&�4�!�]�}�W���Y����\��
P�����
�
�
�
�"�o�N���&����l�N��Uʴ�
�1�0�h�w�/�(���&����U��W�����9�y�u�u�w�}��������X��E��*ڊ�
�
� �g�n�<�(�����ƹF�N�����%�4�d��j�}����&ù��9��h\�*���4�%�4�d��W�W���Y�ƥ�l��h\��U��2�%�3�e�1�l����Oʹ��l��h\��Y���u�u�u�<��8����/���T��Q1�����3�
�c�
�9�?����&��ƹF�N�����!�'�
�u�i�:����I����l ��X�����0� �;�e�]�}�W���Y����V��Y1�H���'�
�
�
�����@����A��E ��Y���u�u�u�4��8����K���T��Q1�����3�
�c�
�'�/����&��ƹF�N�����!�'�
�u�i�:����I����l ��X�����0� �;�f�]�}�W���Y����VF�	��*���
�
�
� �e�d������Ɠ9lǑN��X���=�u� �'�9�}����Yۇ��p5��D�����=�u�!�!�w�<����W���F�V��&���8�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�<�(������F��h=�����3�8�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�0�|�!�2�}�W���Y���F�N��U���%��
�&�w�`����*����l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}����&ù��9��h\�*���&�4�!�4��)�����ƭ�@�������{�x�_�u�w�/�(���&����U��W�����4�!�4�
�#�/�(���&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�P�����3�d�3�
�a���������C9��V�����i�u�%�6�9�)��������F�N��U���0�&�_�u�w�}�W���Y���Z �F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h_��U���6�|�4�1�9�)��������W9��G�����u�u�u�u�w�}�W���Y�����h��*���
� �g�l�6�����&����G��h��U��4�
�:�&��2����B���F�N��U���u�9�<�u��-��������Z��S�����
�
�
�
�"�o�N���&����JO�C��U���u�u�u�u�w�}�W���YӁ��l ��h��*���g�l�4�
�#�/�(���
����l��R�����:�&�
�:�>��L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�e�4�'�<�!���&����C�������%�:�0�&�w�p�W���	�֓�_��h8�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&ù��C��a1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�0�$�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���Yӏ����D�����a�`�u�=�9�W�W���Y���F�N��U���u�%�e�4�'�<�!���&����C��R�����:�&�
�:�>��L���Y���F�N��U���u�9�<�u�6���������F��R ��U���u�u�u�u�w�}�W���Y����lV��[��*���%�#�1�%�2�}�JϮ�I����[��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����R
��V1�����u�&�<�;�'�2����Y��ƹF��h^�����
�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�֓�_��h8�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�-�G���	����l��A��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(������O��_�����u�u�u�u�w�}�W���Y����R
��V1�����u�h�%�e�6�-����s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
��<�(���	����l��PN�����u�'�6�&�y�p�}���Y����^��a1��*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�H����l0��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�4�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���F�N�����3�}�%�&�0�?���PӒ��]FǻN��U���u�u�u�u�w�}�W���&¹��K9��V�����'�2�i�u������&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�l����/����TF��D��U���6�&�{�x�]�}�W���&����e9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�6��(������R��X ��*���g�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��u��������\��h_��U���6�|�4�1�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lW��V��*���#�1�|�u�?�3�}���Y���F�N��U���%�d�8�-��-����DӖ��l��h8�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����c��X
�����1�%�0�u�$�4�Ϯ�����F�=N��U���
�0�<�1�6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*؊�0�<�1�4��1�(������R��X ��*���<�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U���}�%�&�2�5�9�C��Y����l�N��U���u�u�u�u�w�}�WϮ�K����Z	��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*��u�=�;�_�w�}�W���Y���F�N��Uʥ�g��'�:��-����	����[��h\�����1�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���<�1�%�0�w�.����	����@�CךU���
�
�0�<�3�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��1�����
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�o�'�������l��G�����u�u�u�u�w�}�W���Y�����h>�����%�0�u�h�'�o�'�����ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�h����&����l��h��ʴ�&�2�u�'�4�.�Y��s���C9��U��*���%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��C��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z �V�����1�
�b�|�#�8�W���Y���F�N��U���u�u�u�
��8��������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&����_�C��U���u�u�u�u�w�}�W���Y�����h�����4�
�9�
�%�:�K���&ƹ��G��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����Q��h8�����4�&�2�u�%�>���T���F��1�����
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�L����R9��G��U��4�
�:�&��+�E��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�0�4��<�(���P����[��=N��U���u�u�u�u�w�}�W���&����l0��E��I���
�
�0�4��W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X����9�
�:��2��������Q��D��ʥ�:�0�&�u�z�}�WϷ�&����\��X�����2�g�b�4�$�:�(�������A	��D�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���O��_��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�W������F�N��U���u�u�u�<��4�1���5����Z9��P1�B��u��9�
�8�����H¹��T9��UךU���u�u�u�u�w�}����Yۇ��@��U
��D��u�=�;�_�w�}�W���Y���F�N��*����'��:������L�����T�����g�e�_�u�w�}�W���Y���V��^�U���u�u�u�u�2�9���s���F�R ����u�u�0�1�'�2����s���K�V�����'�6�&�{�z�W�W�������@F��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���^�Ƹ�VǻN��U���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o����H�ƭ�WF��CF�����;�!�9�2�4�m�JϹ�	����l ��h��G���4�
�:�0�~�t����s���F�N��U����d��'�0�k�E��Y����cW��h��G���%�}�|�_�w�}�'ށ�&����Q��G��Hʚ�d��3�
�n��F��B���)��h8�����b�}�|�i�w��(�������l��G�U����d��'�0�k�E��Y����cW��h��G���%�}�|�_�w�}�'ށ�&����Q��G��Hʚ�d��3�
�n��F��B���)��h8�����b�}�|�i�w��(�������l��G�U����d��'�0�k�E��Y����cW��h��G���%�}�|�_�w�}�'ށ�&����Q�� G��Hʚ�d��3�
�n��F��B���)��h8�����b�}�|�i�w��(�������l��G�U����d��'�0�k�E��Y����cW��h��G���%�}�|�_�w�}�'ށ�&����Q��^��I����
�
� �e�d����I��ƹF��g_��*���
�b�}�d�w�`�8���/����_��G_��D��u�u��d��/���K����Z�x>��#���
�l�
�d�f�t�}���Y����e9��P1�G��|�i�u������@����U�=N��U���
�
�0�
�`�u�C���Dө��l0��B1�L���}�a�n�u�w��F�������T�G��Hʚ�d��3�
�n��F��P���F��1�����c�g�d�|�k�}�'ށ�&����
_��F�\�ߊu�u��
��8�(��Q���[��g_��*���g�l�%�}�`�f�W���6�ד�l��hX�]��u�h��d��;�(��&���O��N��:����'�2�c�e�l�^��Y����e9��h\�*��d�|�_�u�w��(�������N��N�U���
�
� �g�n�-�_��B���)��h8�����b�}�d�u�j��F�������
9��\�N���u��d��%�:�A��K���F��1�����l�
�d�g�~�W�W���)¹��A��Y�G���i�u��
��(�E���	����]ǻN��%ۊ�
�0�
�b��i�W��6�ד�l ��W�����a�n�u�u��l�!�������T��R��:����3�
�l��l�E���s���|6��a1����g�g�|�i�w��(�������l��X����u��
�
�2��@���N���)��h8�� ��l�%�}�b�l�}�Wϑ�H����V�� \��M���h��d��1��Nց�H����l�N��D���'�2�c�g�e�t�K���)¹��U��W��D��|�_�u�u���(���&���� V�S��%ۊ�
� �g�l�'�u�G��Y����cW��h��*��}�d�u�h��l�!���&����CW�G�U���u�u�u�u�w�}��������G��h=��4���4�0�4�������L�����h��*���
� �g�l�6���������F�N��U���u�u�3�%�9�9�(�������r
��V,�����
�
�0�
�a�}�JϹ�	����l ��h��G���4�
�0� �9�o�}���Y���F�N�����;�1�
�0�:��:�������R ��h�����`�u�h�2�'�;�G���H����P��V�����;�e�_�u�w�}�W���Y���F$��X
�����
���%�6�8����&����T9�� N�U���
�
�
�
��(�E�������G��h]�U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K��D��ʥ�:�0�&�u�z�}�WϮ�����N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W��PӒ��]l�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�����PӇ��N��^�����
� �f�g�'�}�W�������l
��h^��\ʡ�0�_�u�u�w�}�W���Y�ƞ�]��h��*���&�'�2�b�g�a�W����ד�_
��Y�����d�
�g�_�w�}�W���Y���F��Y	��*���
�0�:�
�2��D���DӴ��T��V�����&�3�
�d��o�}���Y���F�N�����9�
�e�'�0�j�G��Y����U�� W��G���u�:�;�:�e�t�}���Y���F�N�����
�0�
�d�w�`��������
9��\����!�u�b�n�w�}�W���Y���F��h��*���0�
�g�u�j�/�������� _��G\�U���u�u�u�u�w�}��������Z9��P1�F��u�0�
�8�e�4����KŹ��l�N��U���u�u�u�&�;�)��������S�
N�����%�<�3�
�f��E�ԜY���F�N��Uʦ�2�7�!�'�0�j�D��Y����U�� W��G��u�:�;�:�a�t�}���Y���F�N�����c�
�0�
�e�}�JϬ�/����Q��G\��Lʱ�"�!�u�l�l�}�W���Y����������u�u�u�;�w�;�}���Y����C��R�����u�x�u�&�>�3�������KǻN�����&�u�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��R���=�;�u�u�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��Q��F���u�=�;�u�w�}�W���Y�����h��3����:�
�l�e�8�G�������S�
N�����
�:�
�:�'�l�(݁�&ù��U��W��F�ߊu�u�u�u�w�}�W�������l ��h"����
�
�
�
�2��F���DӇ��l
��q��9���
�l�g�0�f�l����@Ź��l�N��U���u�u�u�6���2���+����lR��R1�����d�g�i�u�%���������C9��h\��*ڊ�
� �`�g�'�f�W���Y���F�N��������!�%��C���H����lT��R�����9�
�:�
�8�-�Fց�&���� 9��hX�*��_�u�u�u�w�}�W���Y����}"��v<�����a�
�
�
�2��@���DӇ��l
��q��9���
�l�g�0�g�l����O˹��l�N��U���u�u�u�6���2���+����lR��R1�����g�a�i�u�%���������C9��h\��*ۊ�
� �c�a�'�f�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠu�u�x�u�$�4�Ϯ�����F�=N��U���6�&�u�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��R��u�=�;�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1����|�u�=�;�w�}�W���Y���F��{1��*���
�:�%�d��8�(��Y����9��h(��*���%�d�
� �d�e���Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u���(���&����U��X����|�i�u�e�g�m�G��I����V��^�E��e�e�e�n�]�}�W������V��D�����%��
�&�~�2�W���Y����VF��T�����x�u�u�4����������]9��X��U���6�&�u�4������Y����VJ��G1�����1�l�y�2�'�;�G���H����P��V�����u�-�!�:�3�4����I����l�N�����u�u�u�u�4�.�W���:����^F��=N��U���u�u�u�=�9�<�(���
�ד�@��S����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t��������C9��P1����|�|�!�0�]�}�W���Y���F�N������3�8�i�w�-�$�������^9��=N��U���u�u�u�u�w�1����Y���F�N��U���u�%��
�$�}�JϿ�&����GW��D��N���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�=�;�4��	��������[�=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Q����\��h�����u�u�'�
���(ށ�����l��S��\���u�=�;�u�w�}�W���Y���F���;���&�u�h�4��	��������l�N��U���u�u�u�0�$�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����U��UךU���u�u�u�u�w�}�������F�N��Uʢ�0�u�%���)�(���&���l�N��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�2�_ǻ�����W9��Q��E؊�g�h�4�
�8�.�(���&���F��R ךU���u�u�u�u�w�}�W���	����U��S�����
�!�
�&��f�W���Y���F�N�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�c�;���s���F�N��U���0�1�<�n�w�}�W���Y����[��V��!���a�3�8�f�j�}�W���Y���F�N�����
�&�u�h�6��#���J����lT��N��U���u�u�"�0�w�)����D���F�N��U���u�u�4�
��;���YѾ��kD��N��U���0�1�6�&�l�}�Wϻ�Ӗ��P��d��Uʚ�d��3�
�n��F��Y����_	��T1�����}�0�<�0�"�.����Q����c��X
�����2�y�a�|�]�}�W����ד�_
��Y�����d�
�g�i�w�l�W����μ�a��[��B���3�
�e�
�c�`��������_��qG�����w�w�_�u�w�<��������V��h��A���%�u�h�w�u�*����	����F
��Y��*���a�g�%�u�w�-��������lV�R��U��n�_�u�u�z�<�(���Ӈ��Z��G�����u�x�u�u�6���������]9��X��U���6�&�}�%�4�q��������V��c1��F���8�g�u�-�#�2��������9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����:�}�0�<�4�3�(�������l��
N��*���&�
�#�
�~�t�W������F�N��Uʴ�
�:�0�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��Y��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������u�&�<�;�'�2����Y��ƹF��G1�����&�<�;�%�8�}�W�������R��C��Yʴ�
�<�
�&�&��(���&����OǻN�����_�u�u�u�w�;�_ǰ��έ�l��D�����
�u�u�%�$�<�������R��X ��*���<�
�u�u�'�.��������l��h��*���|�!�0�u�w�}�W���Y����C9��[��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����W��D��ʥ�:�0�&�u�z�}�WϿ�&����J9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�
�&��q��������Z9��h]�*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C]�����|�4�1�;�#�u��������l ��^�����u�%�6�;�#�1�F��P����[��=N��U���u�u�u�%�%�<���Y����\��h�����n�u�u�u�w�8����Y���F�N�����4�,�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h_�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�d�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u��������B9��h��*���
�y�2�%�1�m��������
9��h
���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�d�u�j�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����4�
�:�&��2����Y�ƫ�C9��1��D���
�c�
�%�3�3�^���s���V��G�����_�_�u�u�z�<�(���&����U��V�����'�6�&�{�z�W�W���	����l��h_�*���<�;�%�:�w�}����
�έ�l%��Q�����u�0�<�_�w�}�W���Y���F��h��*���
�f�u�h��-��������lW���6���&�}�u�:�9�2�E���s���V��G�����_�_�u�u�z�<�(���&����P��V�����'�6�&�{�z�W�W���	����l��h_�*���<�;�%�:�w�}����
�έ�l%��Q�����u�0�<�_�w�}�W���Y���F��h��*���
�c�u�h��-��������lW���6���&�}�u�:�9�2�D���s���V��G�����_�_�u�u�z�<�(���&����V��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��^�����;�%�:�u�w�/����Q����`9��ZGךU���0�<�_�u�w�}�W���Y���R��^	�����e�i�u�4������Iӂ��]��G��U���6�;�!�9�f�l�L���YӃ����T��N�ߠu�u�x�u�'�.��������R��P �����&�{�x�_�w�}��������lU��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����R
��V1�����9�|�u�u�5�:����Y���F�N��U���&�2�7�1�d�}�J�������]��[����h�%�e�4�'�<�!���&������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^��Y����]��E����_�u�u�x�w�-��������F��D��U���6�&�{�x�]�}�W���
����W�� 1�����
�'�6�o�'�2��������R�������6�0�
��$�l����I�Ƽ�9��O1�����9�|�u�u�5�:����Y���F�N��U���&�2�7�1�c�}�J������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��D���-��4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������T9��R��!���f�3�8�g�w�%��������F9��1��\���u�7�2�;�w�}�W���Y���F��G1�����1�a�`�i�w�u��������\��h_��U���&�2�6�0��	��������F��SN�����-�!�:�1�>�;�(��&�����T�����d�e�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�B���
������T��[���_�u�u�%�$�:����LŹ��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(݁�����l��A�����u�0�<�_�w�}�W���Y���F��h��*���
�c�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lT��R�����
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�A���
������T��[���_�u�u�%�$�:����Oʹ��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(ځ�����l��A�����u�0�<�_�w�}�W���Y���F��h��*���
�l�i�u�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G�����}�%�6�;�#�1����H����lS��R��#���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�N���
������T��[���_�u�u�%�$�:����@����@��h����%�:�0�&�6�����UӖ��l��_��*���#�1�<�
�>�q��������l��A�����<�y�%�g��/����	����l��D��U���
�0�4��6���������l�N�����u�u�u�u�w�}�W�������T9��S1�U��}�%�`�7�#��(�������]9��PN�����:�&�
�:�>��^ϱ�Yۖ��l6��^�����9�
�;�&�0�`��������_	��T1�U���}�
�
�4����������@��
N��*���&�
�:�<��t����	�֓�_��h8�����1�<�
�<�w�}��������\��h^�����4�
�!�'�w�}��������\��h^��N���u�0�1�%�8�8��Զs���K��G1�����0�
��&�f�;�������]F��X�����x�u�u�4��4�(�������@��Q��E���&�2�
�'�4�g��������C9��P1����|�u�u�7�0�3�W���Y����UF��G1�����1�g�|�!�2�}�W���Y���F��G1�����0�
��&�f�;���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�g�3�:�l�����Ƽ�\��D@��X���u�4�
�<��.����&����U��1�����
�'�6�o�'�2��������T9��S1�D�ߊu�u�0�<�]�}�W���Y���R��^	�����d�|�!�0�w�}�W���Y�����D�����
��&�g�1�0�F��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�E������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�f�3�8�e�<����Y����V��C�U���4�
�<�
�$�,�$�������^9��V�����'�6�o�%�8�8�ǿ�&����Q��]����u�0�<�_�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y����C9��P1������&�f�3�:�o�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�n����K���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���a�3�8�f�6�.��������@H�d��Uʴ�
�<�
�&�&��(���&���� 9��D��*���6�o�%�:�2�.��������W9��GךU���0�<�_�u�w�}�W���Q����Z��S
��C���!�0�u�u�w�}�W���YӇ��@��T��*���&�a�3�8�d�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����0�
��&�c�;���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�<����&����	��h_��E���e�g�3�
�b��F��Y����_	��T1�����}�0�<�0�"�.����Q����_��X�����d�
�
�
��(�B���	���O�=N��U���
�!��'��2�(���I����l ��Z�����h� �
�����������G9��h��@���%�}�d�1� �)�W���s���R��[�����:�%�d�
���(���L�ӓ�F���*���<�
�0�!�%�(�����έ�A9��h(��*���%�d�
�
���(���L�ד�O������1�%��9�����A����]ǻN�����!��'��8��N����֓�l ��X�����h�_�u�u�w�}����=����a��Z1�*���
�0�
�b�w�5��������CT��h��*��}�|�h�r�p�}����s���F�V�����:�
�:�%�f��(���&����W��UךU���'�
�!��%�����@�ԓ�lV��h��@���%�u�h�_�w�}�W�������l ��h"����
�
�
�
��(�B���	�ƻ�V�D�����<�'�2�c�b�m�W���H����_��=N��U���u�9��������&�ғ�lV��R	��L��u�u�4�'�;���������
9��R1��F���
�m�
�f�k�}�W���Y����_9��s+��'���'�
�a�0�g�/���Kӑ��]F��R�����<�'�2�c�d�m�W���H����_��=N��U���u�'�
�!��/�;���&�ߓ�l��h\�� ���`�%�n�u�w�<����&����	��h_��G���e�`�3�
�o��D��Y���F���*����'��:��d�G���I�ԓ�F9��1��U���;�}�0�
�:�o��������V�
N��R���9�0�_�u�w�}�W���&����\��X��Dӊ�
�
�
�
�2��G��Y����A��C1�����:�
�l�g�2�m����O¹��Z�=N��U���u�9��������&�Г�lV��R	��B���=�;�}�0��0�(�������N��S��D���0�&�u�u�w�}�WϿ�����u	��{��*���e�0�e�g�1��Bށ�H���F��E1��*���
�:�%�d���(ށ�&����
P��N�U���u�u�u�4�%�1�(���&����lW��1��D���
�`�
�g� �8�Wǭ�����9��E��C��e�u�u�d�~�8����Y���F��E�����'��:�
�n�o��������^��N�����9�
�:�
�8�-�Fց�&����9��hX�*��i�u�u�u�w�}��������A9��X��L���0�d�3�
�b��Eϩ�����V
��Z��*���
�m�}�|�j�z�P������F�N���������2�0�Cہ�&¹��T9��UךU���'�
�!��%�����@�ԓ�lW��h��C���%�u�h�_�w�}�W�������v>��e����
�
�
�0��n�W����ο�_9��G\��*���
�l�}�|�j�z�P������F�N�����9�
�:�
�8�-�Fց�&����9��hX�*��_�u�u�'��)�1���5����_��h��*ފ� �c�b�%�w�`�}���Y���P
��y*��4���0�8�a�
������M�ƻ�V�D�����<�'�2�c�b�m�W���H����_��=N��U���u�'�
�!��/�;���&�ߓ�l��h��@���%�n�u�u�6�/��������\��1�����`�3�
�g��n�K���Y���F��[1��1����!�'�
�a�8�F���������YN�����8�g�<�'�0�k�D��Y���O��[�����u�u�u�'��)�1���5����_��h��*ފ� �c�b�%�l�}�Wϼ�����l��B1�C���u�h�}�0��/�(���&����lR��h����
�l�1�8�%�<�(�������U��^��G��u�u�7�8�%�8��������l ��W�����h�}�
�l�3�0����&����U�� V��Gʴ�1�;�2�&�4�3��������9��UךU���4�'�
� �c�l����D�θ�C9��h��*��u�;�u�8��i����&����CT�=N��U���0�0�
�0�8����O����[�N��U����;�0�
�;��������� V��_��]���'�
� �a�f�-�_���D����F��D��U���u�u��;�2���������A�� ]����u�-�!�:�3�4����I����Z�_�����u�<�
�<��/�;���&����T9�� N�����:�&�
�#��t����Y���9F���*����'��:��k�!���&����CU�
NךU���u�u�-�
�8�8����&����_��u��3���&�'�2�c�e�*����
����^��^1��*��
�g�e�u�w�l�^ϻ�
��ƹF�N�����'�4�
�&�>�3����Kù��lǻN��Xʲ�%�3�e�3�f�;�(��&����VF��D��U���6�&�{�x�]�}�W���&����U9��Q��Cӊ�%�6�
�&�>�3����Y�Ƽ�\��DF��*���
�&�$���)�(���&����C9��N��*���
�1�
�f�w�-��������`2��C\�����|�u�u�7�0�3�W���Y����UF������!�9�2�6�f�`�����ƭ�WF������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�2�_���
����W��G�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�^������F�N��U���2�%�3�e�1�l����Oʹ��l��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�2�'�;�G���H����P��V����u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��ƓF�P�����3�d�3�
�a��������F��G1��E���d�3�
�c��-��������@��C1���ߊu�u�'�
���(ށ�����l��V������i�u�
��1����&����Z��N�����3�e�3�d�1��Aց�����R9��aN�U���
�0�4��>����Y����A��h^��*ۊ� �g�l�<��<�(݁�Y����lW��V��*���&�2�_�u�w���������\��1��*��
�g�i�u�#�����&����\��Y�����<�
�<��%�����&����S��E�����;�1�4�
�8�.�(���&���9F� ��*���
� �a�f�'�}�J�������G9��P1�Fʴ�1�!�%�`�����N����l�N�����6�;�!�<�1��Oׁ�K�����1�����
�c�
�g�8�}��������G9��Q��Mي�g�n�u�u�8��(�������Z��Q��Gڊ�f�i�u�u�w�}�Wϸ�	����V9��E��#���%�4�0�4���(���&����D��F�����%�<�3�
�f��E��Y���O��[�����u�u�u�-��2��������~'��_������g�'�2�a�o�}���Y���C9��V�����4�
�9�
�9�.�Ͽ�
����C��R��U���u�u�%�e�6�-��������W9��h��*���<�;�%�:�w�}����
�μ�9��G��#���
�9�y�%�g�<����/����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u������&����l��G�����_�u�u�u�w�}�W���&����R9��V�����;�&�2�i�w��(�������R��[
�U���u�u�0�&�w�}�W���Y�����h�����
�%�#�1�>�����DӖ��l��_��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lV��[��*���;�&�2�4�$�:�W�������K��N�����4�%�4��>�����
����l��TN����0�&�%�e�6�-����Y����R
��V1�����y�%�e�4�'�<�!���&����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�e�4�%�4��<�(���P�Ƹ�V�N��U���u�u�%�e�6�-��������TF���*���=�
�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�9�=���������C9��V�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}���&����\�
N��*���0�!�'�
����������c9��E��C��_�u�u�x�w��B�������R��[
�����;�%�:�0�$�}�Z���YӖ��9��T��*���#�1�4�&�0�����CӖ��P�������4�
�<�
�$�,�$�������^9�������1�<�3�
�g��E�ԜY�Ʈ�T��N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!��.�(�������\�R�����
�
� �f�e�-�W���	����@��A_��\���u�=�;�_�w�}�W���Y�Ƽ�S��R�����
�9�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�S��R�����
�9�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�6��(�������]9��PN�����u�'�6�&�y�p�}���Y����^��a1��*���
�;�&�2�6�.���������T��]���
�4�
�
�'�+����&¹��K9��V�����'�2�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�H����l0��G1�����!�0�u�u�w�}�W���YӖ��l��h8�����1�<�
�<�w�`��������l��A�����u�u�u�9�2�W�W���Y���F��1�����4�
�9�
�9�.���Y����^��a1��*���
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����^��a1��*���u�&�<�;�'�2����Y��ƹF��h_�����
�;�&�2�6�.���������T��]���
�4�
�y�'�l����/����TJ��h_�����
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l��h8�����1�|�!�0�w�}�W���Y�����h��*���;�&�2�i�w��(���&��ƹF�N�����_�u�u�u�w�}�W���&����e9��h��U��%�d�8�-��-���Y���F��Y
�����u�u�0�1�'�2����s���F���*���<�1�4�
�;�����Ӈ��Z��G�����u�x�u�u�'�o�'�������l��h�����4�&�2�
�%�>�MϮ�������h>�����4�
�9�y�'�o�'�������l��h���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�o�'�������l��G�����_�u�u�u�w�}�W���&����\��G1�����
�<�u�h�'�o�'�������l��d��U���u�0�&�u�w�}�W���Y����lT��R�����
�9�
�;�$�:�K���&����A��h�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ԓ�V��S1��*���u�&�<�;�'�2����Y��ƹF��h\�����1�<�
�<��.����	����	F��X��¥�g��'�:�{�-�E�������C��N��G���'�:�
�%�!�9�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h>�����4�
�9�|�w�5��ԜY���F�N��G���'�:�
�;�$�:�K���&����A��d��U���u�0�&�u�w�}�W���Y����lT��R�����
�<�u�h�'�o�'�������V��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʥ�f�
�
�
�"�i�E���Y���P��N1��*���
�g�4�1��3�ށ�����V��R	��F���_�u�u�
�n�9��������Z9��hZ�*��i�u�1�9�#�9����
����S��G]��ʦ�2�7�!�'�0�j�D��Y����lU��S�����
�
�:�
��(�B���	���N��W�����2�;�<�<�1��@ׁ�KӞ����T�����d�d�n�u�w�-�C���-����T9��N�U���
�!��'��2�(���K����lP��R	��E��_�u�u�x�'�i�"�������V9��V�����&�<�;�%�8�8����T�����h;�����2�0�e�4��1�(�������A	��N�����&�4�
�0�w�-��������`2��C]�����y�0�<�6�9��(���J�ԓ�OǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���J����lT�V �����}�-�!�:�3�4����I����[��G1�����9�d�e�|�~�)����Y���F�N��*ފ�
�<�<�2�2�m���������T�����2�6�d�_�w�}�W������F�N��U���%�a� ��:�3�(���&����_�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}���YӖ��l3��^�����d�i�u�'��)�1���5����_��h��*���
�d�n�_�w�}�ZϮ�M����Z��P1��D���
�9�u�&�>�3�������KǻN��*ފ�
�<�<�2�2�l��������@��h����%�:�0�&�6�����	����l��F1��*���
�&�
�y�2�4����&����lU��h����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GU��D��\ʴ�1�;�!�}�/�)�������� V��G\��U���6�;�!�9�f�m�^�������9F�N��U���u�
�
�
�>�4����H����E
��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�%�c��#�������9��h��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ߊ�0�4��4��1�(���
����@��YN�����&�u�x�u�w�-�B�������R��[
�����2�4�&�2��/���	����@��h[������4�
�9�{�-�B�������R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�B�������R��[
��U���;�_�u�u�w�}�W���&ƹ��G��h�����<�
�<�u�j�-�B�������R��[
�U���u�u�0�&�w�}�W���Y�����h�����4�
�9�
�9�.���Y����Q��h8�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l��V1�����<�u�&�<�9�-����
���9F���*���4��<�
�>���������PF��G�����%�`�7�!��q��������e9��R	����7�!�
�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h[������4�
�9�~�}����s���F�N�����7�!�
�
�9�.���Y����Q��h8�U���u�u�0�&�w�}�W���Y�����h�����<�
�<�u�j�-�B�������C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���%�c���:�3�(���Y����_9��s+��'���'�
�a�0�g�/���K��ƹF�N��C����8�;�
������Ӈ��Z��G�����u�x�u�u�'�k�!�������V9��V�����&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�D������V��T��*��� �f�g�%�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�f�3�8�e�}��������K��X �����
�e�
�g�j�<�(���
����9��G�����u�u�u�u�w�}�WϮ�O����Z��P1��E���
�9�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��c�����
�
�%�#�3�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠu�u�%�c��	����&����[��[1��1����!�'�
�c�8�F�������lǻN��Xʥ�c���8�9��(ށ�	������^	�����0�&�u�x�w�}����/����Z��R1�����9�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���J����lT�R�����
�
� �f�e�-�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�f�1�0�E����Ƣ�GN��O�����<�3�
�e��o�JϿ�&����G9��1�\���!�0�u�u�w�}�W���YӖ��l0��^�����d�4�
�9�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��1��!���;�
�
�
�'�+���Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�'�e� �������V9��S��������!�%��A���I����lW��dךU���x�%�m��#�0����&ù��l�������%�:�0�&�w�p�W���	�ޓ�l��^ �����4�
�9�
�$�4��������C��R�����0�u�%�&�0�>����-����l ��h\����6�;�
�
�"�n�E���P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�n����K�ƭ�WF��CF�����:�1�<�3��m�(��DӇ��P	��C1��D��|�|�!�0�w�}�W���Y�����h9�����2�0�e�4��1�W������]��[����_�u�u�u�w�1��ԜY���F�N��M���!�8�;�
���������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}����.����Z��R1�I���9�����)����O����l��h\�N�ߊu�u�x�%�o�
��������9��h��U���<�;�%�:�2�.�W��Y����l^��h�����0�d�4�
�;���������PF��G�����4�
�0�u�'�.��������l��h��*���0�<�6�;�����K����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������F��SN�����-�!�:�1�>�;�(��&�����T�����d�e�|�|�#�8�W���Y���F���*���<�<�2�0�f�<�(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʥ�m��!�8�9��(ށ�	����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�W���	����F
��Y��*���a�g�%�u�j�/�!���&����CT�N�����u�e�n�u�w�-�!���&����^��^1��*��
�f�i�u�w�}�W���	����9��h��A���%�u�=�;��/����&����]	��^1��*��
�g�e�u�w�l�^ϻ�
��ƹF�N�����;�!�9�f���1���?���F��a��*���3�
�f�
�e�a�W���&����P9��T��]���<�;�1�%��1�(�������V�N�����0�}�8�
�d�4����K˹��O��N�����9�
�
� �b�m����D���F�N��*���&�
�#�g�g�*��������A��B1�F���}�|�h�r�p�}����s���F�G1��؊�d�3�
�f��o�}���Y����_T��h��@���%�u�h�_�w�}�W���&����lT��h��*��� �`�g�%�w�5��������V9��Q��E܊�g�e�u�u�f�t����Y���F������<�3�
�g��n�}���Y����@��Y1�����g�
�g�i�w�/��������lQ����U���!�'�2�b�b�f�W�������F9��1��U��3�%�9�
�8�����HŹ��U��\��F�ߊu�u�
�
�"�o�N���Y����cW��h��*��}�g�x�d�3�*����P���F��a1��*��
�g�i�u�#�����&����\��R�� �&�2�0�}�#�����&����\��^	��§��3�
�b��m�W�������A��H��#���
�b�
�d�~�q�A���B�����B1�A���u�h�w�w� �8�WǪ�	���� Q��G_��U���6�;�!�9�e��^ϻ�
���]ǻN��*���
�
� �f�a�-�W��Q����R��B1�M���u�'�'�3��j�(��B�����h��G���3�
�g�
�e�a�W��Y����N��h��3����:�
�
�2��B���Y����\��h��*���0�&�u�e�l�}�Wϭ�����l��B1�A���u�h�w�w� �8�WǷ�&����\��X�����2�g�b�h�6�����&����O��[��W���_�u�u�<�9�4�(���&����lR��h�I���&�2�7�!�%�:�@������C9��Y�����d�n�u�u�#�-�B܁�&����^��N�U���
�:�<�
�2�)�Ǭ�
����F��P ��]���4�&�2�
��(�C���	���O�=N��U���
�a�<�3��i�(��E����^��1��*��
�f�-�'�6�����&����O��N�����`�
�
� �c�j����D�μ� ^��h�� ��g�%�u�:�w�-��������lW�=N��U���
�a�3�
�o��D��Y����U�� W��G��u�:�;�:�e�t�}���Y����S��B1�B���u�h�%��;��F���&����CT�N�����u�d�n�u�w�)����&����CW�
N��#���
�b�
�g�e�}�W�������V�=N��U���-� �,� ��(��������U��X��G��u�!�
�:�>�����ۓ��Z��SF��G���'�:�
�;�$�:�W�������V��h8��G���3�
�g�
�d�t�}���Y����E]�