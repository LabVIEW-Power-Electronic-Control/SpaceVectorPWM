-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�e������(���
����GF�N�����9�u�u����;���:���F��h��U���������}���Y����G��T��;ʆ�����]�}�W�������	F��cN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�%�<���6����g"��x)��N���u�<�
�%�%�8���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF��Y1�����
�u�u����;���:����g)��]����!�u�|�_�w�}��������G9��N��U���
���
��	�%���Hӂ��]��G�U���<�
�%�'�2�)�E��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����E�����u�u� �u���8���&����|4�_�����:�e�n�u�w�<�(�������\��b:��!�����
����_������\F��d��Uʴ�
�0� �;�e�g�8���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƭ�l��B��F��������4���:����U��S�����|�_�u�u�'�/����&����|3��d:��9�������w�n�W������]ǻN�����!�'�
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W�������\��yN��1�����|�_�9�f�}������P��RN�����:�u��`�`���������@FǻN�����4�!�4�
�8�.�(�������	F��s1��2���o�u�d�n�w�}��������R��X ��*���<�
�u�u���8���Y���A��N�����!�;�u�%���ށ�
����	F��s1��2������u�b�9� ���Y���F�^�D��u�u�6�;�#�3�W���*����9��Z1�Oʆ�������8���Lӂ��]��G��H���e�e�e�n�w�}��������R��c1��F���8�g�o����0���/����aF�
�����e�u�h�w�g�l�G��Y����\��V ������&�a�3�:�n�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���I����]ǻN�����4�!�4�
��.�B������5��h"��<������}�w�2����I����D��^�W�ߊu�u�:�&�6�)����-����l ��h[��U���
���
��	�%���Y����G	�N�U��e�e�w�_�w�}��������C9��Y����
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�e�w�]�}�W���
������T�����d�d�o����0���/����aF�
�����e�u�h�w�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�l�U�ԜY�Ư�]��Y�����;�!�9�d�g�g�$���5����l0��c!��]���:�;�:�e�w�`�U���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)����I����g"��x)��*�����}�u�8�3���Y���V�=N��U���&�4�!�4��2��������	F��s1��2������u�f�9� ���Y���F�L�U���6�;�!�;�w�-��������lW�=��*����
����u�W������F��L�W�ߊu�u�:�&�6�)��������_��h]��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��_�D��n�u�u�6�9�)����	����@��A]��F���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�D��e�w�_�u�w�2����Ӈ��P	��C1��F؊��o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��d�d�e�n�w�}��������R��X ��*���f�e�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�n�w�}��������R��X ��*���g�a�f�o���;���:����g)��_����!�u�|�o�w�m�G��H����D��N�����!�;�u�%�4�3����H¹�� F��d:��9�������w�l�W������F��L�E��d�e�d�n�w�}��������R��X ��*���g��o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�d�l�}�WϽ�����GF��h�����#�d�e�o���;���:����g)��_����!�u�|�o�w�m�G��I����]ǻN�����4�!�4�
�8�.�(���K����\��c*��:���
�����l��������\�_�D��d�d�e�n�w�}��������R��X ��*���g�f�u�u���8���&����|4�_�����:�e�u�h�u�m�G��H����]ǻN�����4�!�4�
�8�.�(���&����`2��{!��6�����u�`�3�*����P���V��^�N���u�6�;�!�9�}��������EP��N�&���������W������\F��T��W��d�e�n�u�w�>�����ƭ�l��D�����e�o�����4���:����S��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
����T��T��!�����
����_������\F��T��W��e�e�e�e�g�f�W�������R��V�����
�#�g�f�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����W��UךU���:�&�4�!�6�����&����F��d:��9�������w�k��������\�^�E��w�_�u�u�8�.��������]��[�*������o���;���:����g)��]����!�u�|�o�w�l�F��H����W��_�D��d�d�d�d�f�f�W�������R��V�����
�#�g���g�$���5����l0��c!��]��1�"�!�u�~�g�W��H����W��L�U���6�;�!�;�w�-��������9��q(��3�����u�u���8���&����|4�]�����:�e�u�h�u�l�F��H����W��_�D��d�d�d�d�f�l�F��H����W��_�D��u�u�6�;�#�3�W�������l
��1��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�D��w�_�u�u�8�.��������]��[�*��o������!���6���F��@ ��U���o�u�e�e�g�l�G��[���F��Y�����%�6�;�!�;�l�(��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��_�E��n�_�u�u�>�3�Ͽ�&����@�=��*����
����u�W������F��L�E��w�_�u�u�#�/����Y����V��S��U���!�<�2�_�w�}��������U��R �����u�3�4�
��;���
����_F��L�����_�u�u�<�9�1��������V��c1��D���8�e�o����0���s���@��V�����2�7�1�g�w�}�8���8��ƹF��^	��ʴ�
�<�
�&�&��(���&����F��d:��9����_�u�u�>�3�Ͽ�&����Q��V��U�����n�u�w�.����Y����U��\��D��������4���Y����W	��C��\�ߊu�u�<�;�;�;�(�������^9��h��*��a�o�����4���:����U��S�����|�_�u�u�>�3�Ϸ�&����\��X��Dۊ� �g�e�%�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������9��h(��*���%�d�
�0��l�E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V�����&�$��
�#�����Y�Ɵ�w9��p'�����u�<�;�9�6���������\��x!��4��u�u�&�2�6�}��������lT��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2���������Q�=��*����
����u�W������]ǻN�����9�0�<�6�9����M����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�g�1��Bׁ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�
�0��l�B��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��Q=��8���,� �
�f�1��Fׁ�K����g"��x)��*�����}�d�3�*����P���F��P ��U���-� ���#�o�(���&����\��c*��:���
�����l��������l�N�����u�&�0�
�2��F��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*���
�&�$���)�(���&����`2��{!��6�ߊu�u�<�;�;�<�(���&����
R�,��9���n�u�u�&�0�<�W���&�Փ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������_��N��1��������}�B�������V�=N��U���;�9�!�%�f����K����	F��s1��2������u�g�9� ���Y����F�D�����8�
�l�'�0�l�N���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��(�����a�
�g�o���;���:����g)��_����!�u�|�_�w�}����Ӡ��A��\�U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_�������V�=N��U���;�9�!�%�e�����K���5��h"��<������}�w�2����I��ƹF��^	��ʼ�8�b�3�
�`��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��^��B���2�d�d�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lP��Q��LҊ�f�o�����4���:����S��X����n�u�u�&�0�<�W���&�֓�V��\�Oʆ�������8���Lӂ��]��G�U���&�2�4�u��<�E�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�
�6�o�A�������
F��d:��9�������w�n�W������]ǻN�����9�4�
�<��.����&����U��N�&������_�w�}����Ӈ��@��U
��D��o�����W�W���������D�����'�2�d�f�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������l��h_�E��������4���Y����\��XN�N���u�&�2�4�w�8����&����@9��hW�*��o������!���6�����Y��E��u�u�&�2�6�}��������A	��E��D��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1�%���¹��_9��R��*���m�3�
�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��Y	��*���
�;�&�g�>�l�(���&����\��c*��:���
�����}�������9F������4�'�9�
�8�����Hʹ��V9��1��*��c�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Z��D��&���!�
�&�
�w�}�#���6����9F������4�
�<�
�3��D���Y����v'��=N��U���;�9�4�'�;���������
9��R1��F���
�e�e�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����R��[�����:�%�d�
���(ځ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�'��)�1���5����_��h��*ۊ� �d�m�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��3����:�
�l�e�8�F�������
^��N�&���������W��Y����G	�UךU���<�;�9�4�%�1�(���&����lW��1��D���3�
�d�g�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h'��0����0�8�a���(���&����	F��s1��2������u�d�}�������9F������6�
��������Mǹ��9��P1�C��������4���Y����W	��C��\�ߊu�u�<�;�;�<����&����	��h_��G���e�c�'�2�f�e�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�����'��:�
�n�o��������V�=��*����
����u�FϺ�����O��N�����4�u�9����%�������l��h��*��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���0����r4��R��A܊�
�
�0�
�n�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��3����:�
�
�2��G���Y����)��t1��6���u�d�1�"�#�}�^�ԜY�ƿ�T���������!�g��(�E���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�
���,�"��D���&����CW�=��*����
����u�FϺ�����O��N�����4�u�'�
�"�o�E���Y�Ɵ�w9��p'��#����u�c�u�8�3���B�����Y�����&�2�
� �e�h����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����%�
� �g�e�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��S1�����
� �g�`�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��R	��*���f�m�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ʃ�C9��G1�����g�
�a�o���;���:����g)��_����!�u�|�_�w�}����Ӓ��lR��Q��D؊�d�o�����4���:����P��S�����|�_�u�u�>�3�Ϫ�	����F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��n����NŹ��\��c*��:���
�����l��������l�N�����u�8�
�l�1��Oׁ�H����g"��x)��*�����}�u�8�3���B�����Y�����f�
� �f�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h�����l�
�g�o���;���:����g)��[�����:�e�n�u�w�.����Y����^��B1�C���u�u��
���(���-���T��X����n�u�u�&�0�<�W�������lW��Q��Dي�d�o�����4���:����S��S�����|�_�u�u�>�3�ϳ�����l ��_�����u��
����2���+������Y��E��u�u�&�2�6�}����I����U��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�o�(���M�ӓ�F��d:��9�������w�l�W������]ǻN�����9��
�
�"�i�G���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y������3�
�g��n�Mύ�=����z%��r-��'���f�1�"�!�w�t�}���Y����R
��Z��@���
�c�
�a�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��h��A���%�u�u����>���<����N��
�����e�n�u�u�$�:����K�ԓ�R��Q��A݊�d�o�����4���:����U��S�����|�_�u�u�>�3�Ϸ�����lR��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��A���&����CT�=��*����
����u�FϺ�����O��N�����4�u�8�
�`�;�(��&���5��h"��<������}�d�9� ���Y����F�D�����8�
�m�3��d�(��Cӵ��l*��~-��0����}�f�1� �)�W���s���@��V�����a�3�
�`��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���`�d�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƿ�\��R��*���`�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��@���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l��C1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������9��h[�*��o������!���6�����Y��E��u�u�&�2�6�}����N����U��G]��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�k�(���L�ߓ�F��d:��9�������w�h�W������]ǻN�����9�!�%�c��(�B���	����`2��{!��6�����u�`�w�2����I��ƹF��^	��ʡ�%�c�
� �b�e����Y����)��t1��6���u�`�u�:�9�2�G��Y����Z��[N��'���9�
�
� �b�i����Y����)��t1��6���u�`�u�:�9�2�G��Y����Z��[N����
� �`�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������V��A���
�d�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������^��1��*��
�d�o����0���/����aF�
�����e�n�u�u�$�:����&����P��N�&���������W������\F��d��Uʦ�2�4�u�
�����J����	F��s1��2������u�g�9� ���Y����F�D�����7�3�
�a��n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h�����d�3�
�l��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���c�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�e��h[�� ��l�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Q��B1�@���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Oƹ��lS��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2���������9��T��!�����
����_�������V�=N��U���;�9�!�%�1��Cށ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�e�3��i�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�
� �c�n�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��D�����a�1�8�'�6����H����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�d��(�A���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʦ�:�0�0�2�����J����	F��s1��2������u�d�}�������9F������!�%�f�
�"�k�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����3�
�m�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������
9��hY�*��o������!���6�����Y��E��u�u�&�2�6�}��������U��[��D��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����P��N�&���������W��Y����G	�UךU���<�;�9�!�'�i�(���N�֓�F��d:��9�������w�h�W������]ǻN�����9�9�
� �`�k����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���b�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ�� T��B1�E���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����N¹��lQ��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��C���&����CT�=��*����
����u�W������]ǻN�����9�'�#�
�"�j�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����6�&�
� �a�i����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N����
� �b�m�'�}�W���&����p9��t:��U���u�:�;�:�g�f�W���
����_F��Y	��*���
� �b�g�'�}�W���&����p9��t:��U���u�:�;�:�g�f�W���
����_F��a1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������]��h�� ��g�%�u�u���8���&����|4�N�����u�|�_�u�w�4����+����9��[1����� �b�a�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������R��1�����0�
�
�
�"�e�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����d�4�9�:�2��(���N�Г�F��d:��9�������w�m��������l�N�����u�8�
�c�1��E߁�K����g"��x)��*�����}�u�8�3���B�����Y��'���0�
�9�
�2�2�(���A�Г�F��d:��9�������w�m��������l�N�����u�4�2�d�6�1����
�ד�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Cہ�����l^��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��O���&����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�n����O����\��c*��:���
�����}�������9F������&�9�!�%�c�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʺ�
�:�1�f�>�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʇ�;�0�
�9��3����&����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�h����Nǹ��\��c*��:���
�����}�������9F������%�l�
�
�"�e�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V��*���<�3�
�f��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�l�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����P��N1�����
�b�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�g�<�3��e�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
�9�
�0�8��(�������l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�o�(���@�ӓ�F��d:��9�������w�m��������l�N�����u�8�f�
�"�d�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�g�
� �n�m����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���3�
�g�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��M���
�f�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�CU��Q��@؊�g�o�����4���:����V��X����n�u�u�&�0�<�W�������D9��hW�*��o������!���6�����Y��E��u�u�&�2�6�}�(�������T��^1��*���
�g�o����0���/����aF�
�����e�n�u�u�$�:��������_	��Y�����c�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����l��X�����;�!�3�
�`��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��U�����<�<�;�!�1��Aׁ�K����g"��x)��*�����}�u�8�3���B�����Y�����`�
� �l�d�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E����� �l�e�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���d�e�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G]�����e�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӗ��R
��_�� ��� �l�c�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����@��C��E���
�l�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������9��!��*���9�6�9��1��G���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʠ�
����#���������l ��^�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������A9��X��L���0�e�3�
�g�d����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����
�:�
�:�'�l�(߁�&ù��U��]�����u��
����2���+������Y��E��u�u�&�2�6�}��������l*��G1�*؊�
�
� �d�c��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*����'��:��d�E���I�ԓ�F9��]��F��������4���Y����W	��C��\�ߊu�u�<�;�;�<����&����	��h_��E���d�3�
�e�d�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�f��(���&����lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���?����\	��W��*���
�
� �d�g��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��	��*���g�g�6�u�w�	�(���0��ƹF��^	��ʴ�
�0� �;�g�-����Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�D�����%�'�!�'������Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������4�
�0� �9�o����Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����u�%�'�!�%��(�������g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����9�4�
�0�"�3�C�������`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����4�u�%�'�#�/�(ځ����5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���;�9�4�
��;���*����|!��h8��!���}�u�:�;�8�m�L�ԜY�Ư�^��R �������
��0�������]��1�����1�%��_�w�}�������F�N��<���u����l�}�W���YӨ��l5��p+��U�����n�u�w�}�WϺ�ù��w2��N��!����_�u�u�w�}����.����\��y:��0��u�u�u�u�3�(�(���-����z(��p+��\�ߊu�u�:�!��}�W���Yӂ��F��~ ��!�����
����_������\F��d��U���u�1�;�u�w��$���5����l0��c!��]��1�"�!�u�~�W�W���Y�ƨ�F�!��U���
���
��	�%���Hӂ��]��G��N���u�0�1�6�:�2����s���F��Z�����8�e�����(���������\��U���u�u�2�;�%�>�_���Y���/��N��!����_�u�u�w�}�"���-����	F��c+��'�ߊu�u�u�u�>�m� ���1����}2��r<�U���u�u�1� ���#���Y����t#��UךU���:�!�}�u�w�}�WϽ�����}F��s1��2���_�u�u�u�w�8����Y����g"��x)��N���u�u�u�1�9�}�W���*����|!��h8��!���}�f�1�"�#�}�^�ԜY���F��T��;ʆ�����]�}�W���Y����\��b:��!�����
����_������\F��G�U���0�1�6�8�8�8��Զs���P	��X ��ʸ�e���������&�Ԣ�lP��N�����u�0�0�<�w�W�W���Y�ƅ�\��y:��0��u�u�u�u���$���<����}2��r<�U���u�u�1�;���#���Y����t#��=N��U���u�:�!����Mϗ�-����O��N�����u�_�u�u�w�}���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF�N�����o������0���/����aF�N�����u�|�|�_�w�}��������V��=dװ���;�u�u�3�g�;����K������\��*���
�&�
�l�m�>��������vV�� +�����3� �
�g�$�n����K�ד�R��DךU���0�0�<�u�6�}�}���Y���z"�	N����u�u�u� ��	�0���G����F�N�����
���u�i�n�[���Y�����1��1���h�u�g�_�w�}�W�������z"��S�F���u�u�%�'�w�<�W�ԜY���F��Y^��Kʳ�
���,�"��D���&����CV�N��U���1�;�u�k�1��:��� ����U��B1�M���y�u�u�u�w�9����GӀ��K+��c����
� �g�m�'�t�}���YӀ��l��X��C޻�
�g�g� �g�g����������/��4���e�&�!�3��i���&���F��Y��ʸ�%�}�u�u�w�}�>���G����F�N��;������h�w�q�W���Y����Z��`'��=��u�a�_�u�w�}�W�������g.�	N�\���u�%�'�u�6�}�}���Y���P
��
P�����>�_�u�u�w�}����Y����C9��CBךU���u�u�<�e�j�}��������l��=N��U���u�0�h�u�%����K����9F�N��U���!�h�u�'��(�E���	����9F���*���-�
�g�&�a��(��Y�Ư�^��R �������
��-����K����9��N�����'�6�8�%��}�W���Yӯ��X�d��U���u������J���U���F�
��E�����h�u�e�W�W���Y�ƨ�F��~*��U��c�|�u�u�'�/�W���Y���F�N�����k�1�4�&�0����L����9F�N��U���!�h�u�
�$�4����&����CW�=dװ���u�x�u�=�w�(����Y����VF��G1��*���|�:�u�=�w�)��������VH�d��Uʴ�
��3�8�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W�������l ��R������&�d�3�:�m�}���Y���F�R�����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����Y���F�N��U���u�u�u�%������DӇ��}5��D�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����V��Y1�����u�&�<�;�'�2����Y��ƹF��G1�����
�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W�������G��h^�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�����g�u�;�u�8�u��������U��Z��G��4�
�:�&��+�(���P�Ƹ�V�N��U���u�u�u�u�w�}��������lV��E��I���'�
�!��%�����@�ԓ�lV��h��*���n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��h�� ���d�%�0�u�$�4�Ϯ�����F�=N��U���'�!�'�
��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����E�����
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���f�3�8�g�w�3�W���Qۃ��G��S1��*��
�g�h�4��2����¹��O�C��U���u�u�u�u�w�}�W���YӇ��A��E ��*���2�i�u�'��)�1���5����_��h��*���
�b�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��*��� �;�g�%�2�}����Ӗ��P��N����u�%�'�!�%��(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F������'�
�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�f�3�:�o�W���Y������C�����
�f�
�g�j�<�(���
����9��G�����u�u�u�u�w�}�W���Y�����E�����
�'�2�i�w�1�>���!����V��Z��*ڊ�0�
�a�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����0� �;�f�'�8�W�������A	��D�X�ߊu�u�%�'�#�/�(܁�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N�����!�'�
�
�%�:�K���	����@��A]��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�f�1�0�E����Ƣ�GN��O�����3�
�f�
�e�`��������_��G��\ʡ�0�u�u�u�w�}�W���Y���F��G1�����
�
�'�2�k�}����=����a��Z1�*���
�0�
�m�l�}�W���Y���F���U���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9lǻN��Xʴ�
�0� �;�c�-����
������T��[���_�u�u�%�%�)����&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���'�!�'�
��/���Y����\��h��G��_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�d�;���Y����]	�������1�3�
�f��o�JϿ�&����G9��1�\���!�0�u�u�w�}�W���Y���F������'�
�
�'�0�a�W���0����r4��R��A܊�
�
�0�
�d�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���4�
�0� �9�h����Y����T��E�����x�_�u�u�'�/����&ƹ��V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���%�'�!�'������E�ƭ�l��D�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�n����K�ƭ�WF��CF�����:�1�3�
�d��E������]��[��E���|�!�0�u�w�}�W���Y���F�N�����!�'�
�
�%�:�K�������v>��e����
�
�
�0��d�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�<�
�<��/�;���&����T9��N�����u�'�6�&�y�p�}���Y����Z9��E1�����
�0�
�e��.����	����	F��X�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������A��N���ߊu�u�u�u�w�}��������]��[����h�4�
�0�~�)��ԜY���F�N��Uʼ�u�}�%�6�9�)���������D�����
��&�c�1�0�B�������9F�N��U���u�u�u�u�w���������\��h��*��u�h�<�
�>���������l��h_�G�ߊu�u�u�u�w�}�W�������N��h�����:�<�
�u�w�-��������`2��C\�����|�u�=�;�]�}�W���Y���F�N�����<��'��8��(���&����[��G1�����9�g�e�_�w�}�W���Y���F��SN��N���u�u�u�u�w�8�Ϸ�B���F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�C������F��R ךU���u�u�u�u�w�}�E�������F�(�����a�
�g�_�w�}�W���Y���F��Z�����d�d�u�h�>�0�@���&����CT��N��U���u�u�u�u�>�3��������F������3�
�e�
�f�k�W������ O��N��U���u�u�u�u�#�-�Fց�����
S�
N����
� �f�g�'�f�W���Y���F�N�����g�'�2�d�f�}�JϪ�	����U��Z��G�ߊu�u�u�u�w�}�W�������l��h_�E��u�8�
�f�1��Dׁ�H���F�N��U���u�!�%�c��8�(��M���G��^�� ��m�%�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�&�<�;�'�2����Y��ƹF��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G��U���;�u�u�u�w�}�W���YӴ��T��V�����
�
�
�m�%�:�F��Y����R��1�����0�
�
�
�o�;�(��&����F�N��U���u�u�1�9�#�9����
����lW��N�U���0�0�
�0�8����O����9F�N��U���u�u�u�0�$�:��������U��S��*���g�c�3�
�a��D��Y����G	�G�U���u�u�u�u�w�}��������A��\�U��%��9�
��(�A���	��ƹF�N��U���u�u�8�
�n�/���M�����h]�����e�
�g�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dךU���x�4�&�2�w�/����W���F�G�����}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�I�����_�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��h[��\ʡ�0�_�u�u�w�}�W���Y�ƭ�A9��h(��*���%�d�
�
���(���&����[��E�����'��:�
�n�o����L����V��h����u�u�u�u�w�}�W���&����\��X��Dӊ�
�
�
�0��j�W������G9��E1�����l�g�0�d�f�;�(��M����9F�N��U���u�u�u�9���/�������R��h^�����a�u�h�4�%�1�(���&����lW��1��E���3�
�e�e�'�f�W���Y���F�N��������!�%��C���H����lW��R�����9�
�:�
�8�-�Fց�&���� 9��h_�M���n�u�u�u�w�}�W���YӅ��z(��o/�����
�c�0�e�%�:�F��E�ƭ�A9��h(��*���%�d�
�
���(���H����CU��N��U���u�u�u�u�4��9���8����A��1��D���2�d�a�i�w�/�(���?����\	��W��*���
�
� �d�f��D�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�<����Y����V��C�U���%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�|�!�2�W�W���Y���F�N��*���0�!�'�
�g�/���M�����h��G���%�n�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]ǑN��X���&�<�;�%�8�8����T�����T��U´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������W������u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$�������^9����U°�<�6�;�
�"�o�C���Y�ƭ�l��D��ۊ�|�|�!�0�]�}�W���Y���F�Q=��8���,� �
�f�%�:�F��Y����`9��b"��:���g�
� �g�o�-�L���Y���F�N��U���
�8�g�'�0�l�A���Dӕ��l��1��*���
�g�_�u�w�}�W���Y���@��C�����d�`�u�h�$�1��������9��d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԜY�����^	�����0�&�u�x�w�}�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�F�������F�N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!��.�(���PӒ��]l�N��U���u�u�u�<��4�1���5����W��R	��D��i�u��9��2�(���	����U��^��G�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N��ʻ�-�u�!�!�w�<�(������\ ��_�����u�4�=�;�y�p�}���Y����`9��Z1�����
�'�6�o�'�2����Q����G��N��*���3�8�u�%�4�q��������U��Z��G�ߊu�u�0�<�]�}�W���Y������t=�����&�u�u�u�w�}�Wϩ��ƭ�l5��D�����e�h�u�u�w�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R��Y��]���&�4�!�h�6�����&����P9��G�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�����B���F�N��U���u�9�0�u�w�}�W���Y���F���;���&�u�h�4��	��������l�N��U���u�u�u�0�3�4�L���Y���F���ʴ�
��&�g�1�0�F��Y���F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�V��&���8�i�u�%���܁�
����9F�N��U���u�u�u�9�2�}�W���Y���F�N��U����
�&�u�j�<�(���
�ԓ�@��d��U���u�u�u�u�w�8�Ϸ�B���F�N��U���;�4�
��$�n����K���9F�N��U���u�u�u�3��u��������\��h_��U���6�|�4�1�9�)�_�������l ��]�����u�%�6�;�#�1�F��P����[��N��U���u�u�u�u�w�}����*����Z�V��!���d�3�8�e�]�}�W���Y���F�R�����}�%�6�;�#�1����H����C9��N�����-�!�:�1�1��Dہ�K����C9��Y�����e�|�u�=�9�}�W���Y���F�N��U����
�&�u�j�<�(���
�ғ�@��d��U���u�u�u�u�w�8��ԜY���F�N��U���u�4�
��1�0�K���	����@��Q��G�ߊu�u�u�u�w�}�W����ƥ�l�N��U���u�"�0�u�'��(���&���� F�d��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�%��
�$�}�JϿ�&����GS��D��N���u�u�u�u�w�}�Wϻ�
���F�N��U���u�u�u�4������E�ƭ�l5��D�����f�_�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�"�2�}����&����U��N��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�%������DӇ��`2��CX�����n�u�u�u�w�}�W���YӃ��Vl�N��U���u�u�u�u�w�<�(������F��h=�����3�8�a�_�w�}�W���Y���F��SN��N���u�u�u�u�w�*����	����@��Q��@��u�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�-�9���
�����d:��ي�&�
�n�u�w�}�W���Y�����Rd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�c�3�8�b�W�W���Y���F�N��ʼ�n�u�u�u�w�}�Wϩ��ƣ�[��S�U���u�u�u�u�w�}�WϿ�&����@�
N��-����n�u�u�w�}��������9F���U���6�&�n�u�w�}�WϘ�&����@��B1�B���u�h�&�1�;�:��������A��M�����1��
�
�"�i�G���P����]ǑN��3؊�
� �a�e�'�}�J�ԜY���F��h��*��d�"�0�u�#�-�E߁�����l��G��U��|�0�&�u�w�}�W�������9��hZ�*��_�u�u�g�1��Cׁ�K���@��[�����6�:�}�;�>�3�ǿ�&����G9��\��F���x� �&�2�2�u����&���� R��G����u�4�2�d�6�1����&¹��lQ��h�I���!�%�g�3��i�(������^��1��*��
�g�n�u�w�����&����\��h\��*���3�
�d�
�e�a�Wǽ�����l��B1�A���u�;�u�4�0�l��������9��Q��M؊�f�n�u�u��3�ށ�����V��h�� ��g�%�u�h�]�}�W���Y����VW��[�����3�
�d�
�e�*��������]��h�� ��m�%�}�|�j�z�P������F�N�����!�%�`�3��j�(��s���a��R_�����;�&�3�
�f��E��Y۴��T��V�����
�
�
� �o�m�����ƞ�]��h��*���&�d�3�
�c��E��Y����R��1�����'�&�d�3��i�(��E���F��R ������3�
�g��n�JϿ�&����G9��Z��\ʰ�&�u�e�n�w�}�%���¹��_9��E��G���3�
�l�
�d�a�W���Y�����1�����f�
�g�"�2�}��������l��B1�M���}�|�h�r�p�}����s���F�D�����c�3�
�l��n�}���Y����VW��[�����
� �m�c�'�}�J�������l��h�����3�
�a�
�e�%�Ͽ�&����G9��1�N���u��;�0���(���N�ԓ�F���*���<�
�0�!�%�.����������^	��¸�;��3�
�e��D�������V�������1�r�r�s�#�-�Cځ�����l��_��U���;�:�e�|�~�f�W���+����9��[1�����
�
� �m�g�-�W��s���F�e��؊�9�
�;�&�1��Nہ�Kӑ��]F��E1����
�
� �b�e�-�_���D����F��D��U���u�u�'�#��(�@���	��ƹF��V ��G���9�:�0�
�"�j�C���Y���D��_��]���2�g��d�1��O݁�K����l0��B1�M���|�0�&�u�g�f�}���Y����C9��Y�����;�%�:�0�$�}�Z���YӇ��W	��h�����%�:�u�u�%�>����	����A�V�����&�$��
�#�����UӇ��P�V�����&�$��
�#�����UӃ��G��S1��*��
�g�_�u�w�8��ԜY���F��F�����}�%�6�;�#�1����H����C9��V��\ʴ�1�}�%�6�9�)���������D�����
��&�d�1�0�G������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GU��D��\ʴ�1�;�!�}�/�)��������9��S�����;�!�9�d�g�t�^������F�N��U���4�
�:�0�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����S��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C�����9�u�&�<�9�-����
���9F������
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9��=N��U���<�_�u�u�w�}�������R��X ��*���<�
�u�u�'�.����PӇ��N��h�����:�<�
�u�w�-��������`2��C_�����|�|�!�0�w�}�W���Y�����^
��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}���������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����V�������%�:�0�&�w�p�W�������R��V�����'�6�o�%�8�8�ǿ�&���R��^	������
�!�
�$��[ϻ�����W9��h\�*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C]�����|�4�1�;�#�u��������F9��1��U���%�6�;�!�;�l�G���PӒ��]FǻN��U���u�u�%�'�6�$�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������,�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�0� �9�m�����Ƽ�\��D@��X���u�4�
�0�"�3�G���
����C��T�����&�}�%�6�{�<�(���&����l5��D�����g�u�-�!�8�9����Jǹ��F��E1��*���
�:�%�d���(߁�&����S�������'�
�
�'�0�W�W�������F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�������V��T��*���g�a�%�u�w�-��������lV�G�����_�u�u�u�w�}�W�������]9��S�����!��'��8��N����֓�l��h_�N���u�u�u�0�$�}�W���Y���F��G1�����
�u�h�4��8����I����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�'�!�%��W�������A	��D�X�ߊu�u�%�'�#�/�(ށ�
����l��TN����0�&�4�
�2�}��������B9��h��*���
�y�0�<�4�3�(���K�ғ�J��E�����'��:�
�n�o��������V�V�����;�d�%�0�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�f�3�8�e�}��������K��X �����f�
�g�h�6�����&����O�N�����u�u�u�u�w�}��������lW�
N�����
�:�
�:�'�l�(݁�&¹��T9��UךU���u�u�9�0�]�}�W���Y���R��R����i�u�%�'�#�/�(ށ�����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʴ�
�0� �;�e�<����Y����V��C�U���4�
�0� �9�o��������\������}�%�6�y�6�����
����g9��1����u�-�!�:�3�;�(��&���P
��y*��4���0�8�a�
������M����C9��C��*؊�'�2�_�u�w�8��ԜY���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��ي�&�
�|�4�3�3��������]��B1�A���u�u�%�6�9�)����I�����YNךU���u�u�u�u�'�/����&�����~ ��-���!�'�
�a�2�m����H����F�N�����u�u�u�u�w�}�WϿ�&����A��R�����0� �;�g�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����
�u�&�<�9�-����
���9F������'�
�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
�Փ�@��N�����;�
� �g�c�-�[Ͻ�&����k'��C��*���0�d�'�2�f�o�W�������]9��G��\���u�7�2�;�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��Q��G���;�u�:�}�2�4����&���� R��N�����:�&�
�#��t�^������F�N��U���4�
�0� �9�n�K�������v>��e����
�
�
�0��e�L���Y�����RNךU���u�u�u�u�'�/����&�����E�����
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����V��Y1����2�u�'�6�$�s�Z�ԜY�ƭ�l��B��A���&�2�
�'�4�g��������C9��N��*���
�&�$���)�(���&����K��X �����f�
�g�u�;��3���+����^9��h��*���
�f�y�4��8����M����TOǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���J����lT�V �����}�-�!�:�3�;�(��&�����T�����d�e�|�|�#�8�W���Y���F������'�
�u�h�4��9���8����A��1��E���2�d�a�_�w�}�W������F�N��U���4�
�0� �9�i�K���	����F��1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<�(���������^	�����0�&�u�x�w�}��������lS��D�����:�u�u�'�4�.�_�������C9��P1������&�f�3�:�o�W�������l ��]�����6�
��������MŹ��9��P1�A���%�'�!�'������s���Q��Yd��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�����PӇ����F�����;�
� �g�c�-�W���	����@��A_��\���u�=�;�_�w�}�W���Y�ƭ�l��B��@��u�9��������&�Г�lW��R	��L��u�u�u�u�2�.�W���Y���F������'�
�u�h�6������ӓ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���OӇ��Z��G�����u�x�u�u�6���������9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�C��u�4�
�:�$��ށ�Y�ƭ�l%��Q��Aʱ�"�!�u�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���MӇ��Z��G�����u�x�u�u�6���������9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�A��u�4�
�:�$��ށ�Y�ƭ�l%��Q��@ʱ�"�!�u�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���Y����T��E�����x�_�u�u�'�.��������R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��Z��H���%��
�&��}�������F��h�����#�
�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��OϿ�
����C��R��U���u�u�4�
�>�����A����Z��G��U���'�6�&�}�'��(���P�����^ ךU���u�u�u�u�w�}��������lS��S�����:�&�
�#��}�W���:����^N��S�����|�n�u�u�2�9��������9l�N�U���&�2�7�1�`�}����Ӗ��P��N����u�%�&�2�5�9�@ہ�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������Z������!�9�d�d�j�<�(��������Y��G���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�a�6�.��������@H�d��Uʴ�
�<�
�1��i��������\������}�%��
�$�t�W�������9F�N��U���u�u�u�%�$�:����@���N��h�����#�
�u�u�'��(���Q�ƨ�D��]��N���u�0�1�%�8�8��Զs���K��G1�����0�
��&�f�;�������]F��X�����x�u�u�4��4�(�������@��Q��E���&�2�
�'�4�g��������C9��P1����|�u�u�7�0�3�W���Y����UF��G1�����1�g�|�!�2�}�W���Y���F��G1�����0�
��&�f�;���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�g�3�:�l�����Ƽ�\��D@��X���u�4�
�<��.����&����U��1�����
�'�6�o�'�2��������T9��S1�\���u�7�2�;�w�}�W�������C9��P1�����|�!�0�u�w�}�W���Y����C9��P1������&�g�3�:�l�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�o����H���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���f�3�8�g�6�.��������@H�d��Uʴ�
�<�
�&�&��(���&����9��D��*���6�o�%�:�2�.��������W9��d��Uʷ�2�;�u�u�w�}��������T9��S1�\ʡ�0�u�u�u�w�}�W�������T9��R��!���f�3�8�g�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�f�1�0�E��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��A���8�f�4�&�0�}����
���l�N��*���
�&�$���)�(���&����@��h����%�:�0�&�6���������l�N�����u�u�u�u�>�}��������W9��N�����u�u�u�u�w�}��������V��c1��A���8�f�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӇ��@��T��*���&�a�3�8�d�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����
����g9��1����4�&�2�u�%�>���T���F��h��*���$��
�!��.�(ہ�
����l��TN����0�&�4�
�>�����H��ƹF��R	�����u�u�u�3��-��������P�C��U���u�u�u�u�w�<�(���&����l5��D�����a�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������T9��R��!���`�3�8�a�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��Q��@ʴ�&�2�u�'�4�.�Y��s���R��^	������
�!�
�$��(�������A	��N�����&�4�
�<��9�(��P�����^ ךU���u�u�3�}�'�.��������F��R ��U���u�u�u�u�6�����
����g9��1�����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϿ�&����P��h=�����3�8�`�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���4�'�9�
�8�����Hʹ��V9��1��*��l�%�u�h�$�9��������G	��E�����;�<�;�1�6�/��������\��1�����3�
�e�l�'�t�D���B�����h��3����:�
�l�g�8�G���&����l��S��9��� �,� �
�"�)����KŹ��lW��1��]��1�"�!�u�~�W�W�������l ��h"����
�
�
�
�"�l�C܁�K���@��[�����6�:�}�;�>�3�ǿ�����u	��{��*���e�0�e�g�1��G���	�����^	�� �
�f��!�e�����&����lW��1��\��u�u�4�'�;���������
9��R1��D���
�e�c�%�w�`�}���Y���P
��y*��4���0�8�a�
������J�ƻ�V�D�����
�0�
�d�b�m�W���H����_��=N��U���u�'�
�!��/�;���&�ߓ�l��h��D��
�f�_�u�w�/�(���?����\	��W��*���
�
� �d�a��D��Y���F���*����'��:��d�G���I�ԓ�F9��W��Dʢ�0�u�&�9�#�-����H����O�I�\ʰ�&�u�u�u�w�}����7����a4��E��A���e�'�2�d�a�W�W�������l ��h"����
�
�
�
��(�F��&���FǻN��U���9�����)����M����l��h_�U���;�}�0�
�:�o����H����O�I�\ʰ�&�u�u�u�w�}��������A9��X��L���0�e�g�3��m�D���B�����h��3����:�
�l�e�8�G�������Q��N�U���u�u�u�4�%�1�(���&����lW��1��E���3�
�e�l�'�}����Q����G��h��*��`�e�u�u�f�t����Y���F���*����'��:��d�E���I�Г�V��V�U���4�'�9�
�8�����Hʹ��V9��Q��E���%�u�h�_�w�}�W�������v>��e����
�
�
�0��n�W����ο�_9��G1����`�}�|�h�p�z�W������F�N�����
�:�
�:�'�l�(߁�&ù��U��]����u�u�4�'�;���������
9��R1��D���
�e�a�%�w�`�}���Y���R��[�����:�%�d�
���(���H����CT��_��]���
�8�g�'�0�l�A���P���A�R��U���u�u�u�4�%�1�(���&����lW��1��D���2�d�e�_�w�}��������l*��G1�*؊�
�
�
� �f�d�(��E��ƹF�N�����!��'��8��N����ד�F9��]��Gʢ�0�u�&�9�#�-����H����O�I�\ʰ�&�u�u�u�w�}����7����a4��E��A���d�'�2�d�e�W�W�������l ��h"����
�
�
�
��(�F��&���FǻN��U���9�����)����M����l��h_�U���;�}�0�
�:�o����H����O�I�\ʰ�&�u�u�u�w�}��������A9��X��L���0�d�g�3��m�F���B�����h��3����:�
�l�e�8�F�������S��N�U���u�u�u�6���2���+����lR��R1�����d�a�"�0�w�.����	����lW�� F�U���d�|�0�&�w�}�W���YӇ��l
��q��9���
�l�e�0�f�;�(��J����9F���*����'��:��d�E���H�ӓ�F9��\��F��u�u�u�u�w�>�(���<����G��hZ�����'�2�d�a� �8�Wǭ�����9��P1�C���|�h�r�r�w�1��ԜY���F��E1��*���
�:�%�d���(ށ�&����V��G]�U���7�8�'�0�1��O߁�K�����R�����:�
� �l�e�-�W���	����W��E	��*���:�
� �l�c�-�^�ԜY�Ʈ�^��R1�����!�3�
�c��o�K���	����W��E	��*��� �l�b�%�w�3�W�������D9��C1��*��
�g�n�u�w�>����H����F9��1��U��}�0�
�8�f����N����R��C��FҊ� �c�f�%�~�W�W���&����T��B1�@���u�h�3�
������&�Փ�V��Y����u�0�0�0��8��������l��S��U���u�u��;�2���������l��B1�G���u�=�;�}�6�/�(ށ�&����R��F�U���d�|�0�&�w�}�W���YӴ��T��V�����&�g�<�3��d�(��s���V��T��*���g�a�%�u�j��Uϩ�����9��h(��*���%�&�'�2�e�k�JϿ�&����G9��1�U���0�w�w�_�w�}��������U��Z��A��u�'�2��1��Gׁ�H����W	��C��G��u�u�3�
������&�Փ�F9��1��U��3�
�:�0�#�/�(�������R��=N��U���-� ���#�o�(���K�ޓ�F�d��U���u�<�
�%�%�8���������h��G���
�`�
�g�g�}�W��PӃ��VFǻN��U���0�
�8�d�1��B݁�J��ƹF�N�����
�g�
�0�6�.��������@H�d��Uʲ�%�3�
�g��8��������\������}�%�&�4�#�}��������B9��h��*���
�y�4�
�2�}��������B9��h��*���
�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������R��
N��*���&�
�:�<��t�^ϱ�Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\���!�0�u�u�w�}�W���YӁ��l ��\�����h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���&����T��RN�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���T��Q��G؊�e�i�u�!��2����������^�� ���2�0�}�;��/����P����]ǻN��9���
�:�
�:�'�l�(���K�֓�F���*���<�
�0�!�%�(�����Υ�l
��q��9���
�
�0�
�g�t�\ϫ�
����WN��h�����#�
�|�n�w�}����N���� Q��G\��H���w�"�0�u�$�:��������l ��X�����k�&�2�0��-��������9��N�����e�n�u�u�>�0�(���M�ד�F�L�U���;�}�8�
�b�;�(��&�����T�����b�e�u�9�2��U�ԜY�ƥ�V��h��F���%�u�h�1�6�.��������l��=N��U���3�
�f�
�f�a�W���&�ԓ�F9��1��]���u�u�:�;�8�m�L���YӋ��l0��h��A���%�u�h�&�3�1��������AN��D�����%�6�;�!�;�h�(���Tӓ��Z��SF��'���9�
�f�3��l�(��P���F��Y1�����g�
�f�i�w�}�W���YӋ��l0��h��A���%�u�=�;��.��������V�N��R��u�9�0�_�w�}�W���&����_��1��*��
�d�_�u�w�/����@¹��U�� \��G��u�!�%�a��(�@���	�ƭ�WF��A_�� ��e�%�|�_�w�}��������Z9��hV�*��i�u�!�%�c����O����R��E�����g�
�g�n�w�}���&����l^��h�I����;�0�
�;�����&¹��l^��h����0�
� �b�g�-�^�ԜY�Ƽ�
Q��R�����<�3�
�`��o�K�������l ��[�����'�1�9�!�3�'��������R��d��Uʥ�l�
�0�:�0�3��������
Q��G\��H���
�b�1�8�%�<�(�������l��O�����:�&�
�#��t�}���Y����l��B1�G���u�h�}�8��k����Kù����<�����4�9�/�'�$�;�(��&���9F������!�d�
� �c�n����Dӕ��l
��^�����'�'�&�/��3����ے��lW��Q��E܊�f�y�a�|�]�}�W�������l��B1�A���u�h�}�4�����J����R��C��Cي� �`�m�%�~�W�W���&����lW��Z�����m�
�f�i�w�}�W���YӖ��R
��1����g�u�=�;��/����&����]	��Q��CҊ�g�e�u�u�f�t����Y���F������!�9�f�
���1���s���C9��[\��*���`�g�%�u�j�W�W���Y�Ƹ�C9��h��@���%�u�=�;��0�(�������9��^��H��r�u�9�0�]�}�W���Y����V��P�� ���`�%�n�u�w�-�!���&ƹ��lP��h�I���!�
�:�<��8��������]��G1��؊�
� �`�g�'�t�\ϫ�
����WN��G1�*���c�`�%�|�l�}�WϮ�/����9��hX�*��i�u�u�u�w�}��������l ��[�����=�;�}�0��0�Fہ�����R��B1�D���}�|�h�r�p�}����s���F�D�����2�
�
� �c�n���Y����l	��Q��L؊�g�i�u�!��2����������^	��¡�%�`�
� �d�e����Rӓ��Z��SF��*���&�
�#�
�~�f�W���Y����\��T��*���c�`�%�u�j�.��������V��EF�����}�<�;�1�'�.�(���O�֓�O�G����u�%�&�
�"�k�G���Y����G��X	��*���!�'� �&�0�8�_�������V��E�����;�1�4�
�8�.�(���K����]ǻN��U���:�g�6�&��(�A���	�����h�����0�!�'�'�$�'�_�������\��Q��Mӊ�g�y�g�|�]�}�WϮ�
����lP��h�I���!�
�:�<��8��������]��q\�����g�d�u�u�9�4��������]��[�*��|�_�u�u�5�<����&¹��lS��h�I���'�<�<�3��d�(������Q9��h[�*��n�u�u�$��(�B���	���l�N��Uʼ�;�2�'�2�f�e�W����θ�C9��h��@���%�}�|�h�p�z�W������F�N�����
� �`�a�'�f�W�������F9��1��U��&�1�9�2�4�+����Q����G9��P�� ���2�0�}�%�4�3����Lǹ��u ��q(��3���|�!�
�;�2�8�_�������A��H�����`�3�
�b��l�D��Y����G	�G��\�ߊu�u�
� �b�k����D�Υ�^��E��D��u�;�u�8��k����Nù��]ǻN��*���
� �`�f�'�}�J�������l ��V�����'�'�3�
�`��E��Y����V��Q��Cڊ�g�i�u�!�'�j�(���N�ԓ� F��EN��*���&�
�#�
�~�W�W�������lQ��h�I���!�%�c�
�"�j�E���Y����R��X ��*���
�|�_�u�w�8�(���Hù��lP��h�I���!�%�3�
�c��EϿ�Ӓ��lT��Q��Fڊ�g�n�u�u�$�1����H����S��G]��H�ߊu�u�u�u��<�E�������
9�������0�
�8�d��(�A���	����[�I�����u�u�u�u�w�.����	Ĺ��lP��h����u�0�
�8�f���������F9��1��U��}�8�
�g�%�:�F��Y����^��1��*��
�g�n�u�w�.����	¹��lT��h�I���u�u�u�u�>�����������YN�����8�
� �g�a�-�_���D����F��D��U���u�u�<�
�'�/����K���F��[1�����3�
�c�
�e�a�WǪ�	����U��\��Fʺ�u�8�
�a�9�)����LŹ��]ǻN�����8�g�
� �o�e����D�θ�C9��h��M���%�u�;�u�2����&����T��G�U���&�9�!�%�b�;�(��&���FǻN��U���4�2�d�4�;�2����&����P��N�����&�9�!�%�c�;�(��&���F�_��U���0�_�u�u�w�}��������l��=N��U���
�8�g�
�"�e�G���Y���F�N��'���0�
�9�
�2�2�(���A�Г�F��R �����!�%�a�3��k�(��I���W����ߊu�u�u�u��h����&����CT��N�����!�%�b�3��o�(��E����^��1����a�u�:�u�'�>�����ד�]ǻN�����8�g�
� �n�h����D�θ�CU��Q��Fڊ�g�4�1�<�9�:����H����l�N�����%�l�3�
�c��E��Yے��lU��E��D��u�;�u�&�2�����H���9F���*���g�3�
�`��o�K���H�ƻ�V�^"�����'��:�
��8�(��Y�ƭ�l��D��؊�|�0�&�u�g�f�W���
����^��h��L���%�u�h�_�w�}�W���	����@��A]��Eʢ�0�u�!�%�b����J����O�I�\ʰ�&�u�u�u�w�}��������A��\�N���u�&�9�!�'�l����I�ӓ�F�F����
�0�
�d�b�%�Ͽ�&����G9��1�N���u�&�9�!�'�o����I�֓�F�F�����0�3�
�m��o����
����^��h��D��
�g�n�u�w�.����	Ĺ��lP��h�I���u�u�u�u�#�-�Bہ�����l��@��U¡�%�g�
�0��o�E��Y���O��[�����u�u�u�
�6�o�B���&����CT��N�����!�%�
� �a�k����D�θ�C9��h��*��g�-�'�4��2����¹��l�N�����%�3�
�a��o�K���H�ƻ�V�^"�����'��:�
��8�(��Y�ƭ�l��D��؊�|�0�&�u�g�f�W���
����^��R1��*��
�f�i�u�w�}�W�������]��[�*������"�2�}��������lW��F�U���d�|�0�&�w�}�W���YӇ��P	��C1��F؊�n�u�u�&�8�8����&����lR��h�I���u�u�u�u�#�-�Eف�����l��@��U¼�8�
� �a�f�-�_���D����F��D��U���u�u�4�
�8�.�(���K����F�C��G���
�a�
�g�k�}��������l��V �����3�
�g�
�e�f�W�������l ��]�����h�}�0�&�0�?��������F��SN�����%�b�3�
�e��E��Y����^��h��L���%�u�h�}�$�8�(���&����	��D�����b�3�
�g��o�L���YӒ��lW��Q��E܊�f�i�u�4��2����¹��F��G1�*���
�d�e�n�w�}����Hʹ��lU��h�I���d�u�=�;��0�(�������9��S�����;�!�9�c��t����Y���9F���*���3�
�f�
�e�a�W��Y����N��P ��]���'�2�d�e�~�c�����έ�l��D�����e�|�0�&�w�m�L���YӒ��lT��Q��Fߊ�g�i�u�!��2����������^	��´�
�:�&�
�!�o�G���Y����T��(�����d�e�|�n�w�}����K����lU��h�I���d�u�=�;��%�(���&����lU��h�Hʴ�
�:�&�
�!�l�C��Y����D��d��Uʡ�%�g�
� �c�h����D������YN�����;�1��
��(�C���	�����^	��´�
�:�&�
�!�o�D���Y����D��d��Uʡ�%�g�
� �c�j����Dӕ��l
��^�����'�&�<�!�;�;�_���������h[�����`�
�d�y�8�4����ۓ��Z��SF��R���
�
�4�#�;�(��&���K��S�����|�|�|�_�w�}����N����_��G_��Hʦ�1�9�2�6�!�>����������^	���
�
�4�!�1��C؁�H����O��N�����g�
� �a�b�-�W��
����\��h�����&�<�!�'�0�)�����Ρ�]9��Q��Gي�f�y�:�<�#�:�ǫ�
����WN�N�����g�
� �a�f�-�_��Hӂ��]��G��\��u�u�!�%�d����I����[�L�����}�<�;�1������K���F��P ��]���6�;�!�9�f��A�������V�=N��U���
�d�3�
�e��E��Y����_	��T1�����}�;�<�;�3��(���&����F�B �����}�%�6�;�#�1�F݁�?���9F���*���3�
�b�
�e�a�W���&����P9��T��]���<�;�1���(�D���	�����^	��´�
�:�&�
�!�o�1���P���F��G1�*���f�g�%�u�j��Uϩ�����Z��SF����
� �f�c�'�t�Iϭ�����R��X ��*���g�f�|�u�;�8�U���s���G��X�� ���e�%�u�h�u�� ���Yۖ��V��C1�����c�
�g�h�6�����&����lV�R��U��n�u�u�!�'�n�(���O�ӓ�F���*���<�
�0�!�%�/����Q����T�������2�
�
� �b�d����J���9F���*���3�
�g�
�e�a�WǪ�	����U��[��Fʭ�'�4�
�:�$��ށ�P���F��G1�*���b�c�%�u�j��Uϩ�����Z��SF��ۊ� �c�e�%�~�a�����έ�l��D�����f�|�u�9�2��U�ԜY���F��G1�*���!�3�
�f��l�K�������T��A�����0�<�0�&�0�8�_���&�ד�F9��1��\��|�n�_�u�w�0�(�������9��R�����9�2�6�#�4�2�_�������]��Y�����
�4�!�3��e�(��U���l�N����
� �b�e�'�}�Jϭ�����Z��R��¦�<�!�'�2�#�.����Q����e9��hZ�*��y�:�<�!�0�/��������V�N����
� �b�c�'�u�F������\F��G��N���u�!�%�a��(�@���	���D�������<�;�1�%�$����@����Z��^	��´�
�:�&�
�!�o�D���Y����D��d��Uʡ�%�a�
�:��(�O���	���N��G1�*���b�c�%�u�8�}��������EW��UךU���8�
�`�3��j�(��E�ƿ�W9��P�����:�}�0�<�2�(�����μ�@T��V�����l�
�d�y�c�t�}���Y����P��B1�E���u�h�w�w� �8�Wǌ�����e9��Q��M؊�g�h�4�
�8�.�(���M���V
��L�N���u�!�%�a��(�D���	�����P1�����e�
�d�c�w�}�W������]ǻN�����m�3�
�f��o�K���H�ƻ�V�G��*���c�l�%�u�w�-��������9��N�����e�n�u�u�#�-�Cց�����l��S��'���0�
�9�
�9�.�E���H˹��T9��_�����%�6�;�!�;�l�F��Y����^��1��*��
�g�i�u�#�-�Fց�����
S��EN�����9�"�3�
�c��D��Y����^��1��*��
�d�i�u�%�:�!���&����CW�N�Dʱ�"�!�u�|�]�}�W���&�ғ�F9��1��U��8�;��3��o�(��J���F��@ ��U���_�u�u�8��h����O¹��Z�q\��*���a�e�%�}�f�9� ���Y����F�C��@܊� �`�d�%�w�`����K˹��lR��h�F���u�u�:�;�8�m�L���YӒ��lS��Q��Fފ�f�i�u�4�����J����G	��Y�����;�<�;�1�#�-�Cށ�����F9��1��\���:�;�:�!��3����Q����T����*���6�&�
� �b�m����Pӑ��]F��X1�����'� �&�2�2�u����H����G9��h[�*��|�h�e�4�3�)�(�������F��P ��]���
�d�6�&��(�B���	���S�������w�_�u�u�:��O���&����CR�
N��*���f�m�%�}�f�9� ���Y����F�C��@ӊ� �f�m�%�w�`����J����lU��h�C���d�1�"�!�w�t�}���Y����V��B1�M���u�h�_�u�w�}�W�������l
��h]����u�!�%�f��(�D���	����[�I�����u�u�u�u�w�-��������l��=N��U���
�d�3�
�c��F��Y����_	��T1�����}�0�<�0�"�.����Q����V��R	��G��y�a�|�_�w�}����K����S��G\��Hʦ�1�9�2�6�!�>��������_�������1�4�
�:�$�����J����u ��q(��3���:�<�!�2�%�(�������F�C��Cۊ� �`�l�%��l�FϺ�����O�G�U���!�%�c�
�"�h�O���Y���G��\�� ���g�%�u�:�w�-��������9��q(��3�����|�_�w�}����L����^��G]��Hʥ��9�
�
�"�h�E���Q����\��XN�\�ߊu�u�8�
�a�;�(��&���F��a��*ފ� �`�g�%��}�W�������V�=N��U���
�b�3�
�f��D��Y����_T��h��C���%�}�d�1� �)�W��B�����hX�����d�
�f�i�w�2�F���&����CT�N�����u�d�n�u�w�)���&����T��N�U���g�3�
�m��o�F�������W��d��Uʡ�%�3�
�a��o�K�������9��h[�*��4�1�&�9�#�-�(���O�Г�O��N�����&�3�
�f��l�K�������T��A�����0�<�0� �$�:��������C9��Q��Gފ�a�y�g�|�]�}�W����ԃ�G9��h�����
� �d�d��n�K���Y���F��h8��G��
� �
� �n�k�������@��C��G���
�e�e�%��t�J���^�Ʃ�@�N��U���&�9�!�%�g�;�(��&����F�B"��&����!��7�%�>�(�������R��N�U���
�:�<�
�2�)�ǫ�
����WN��h>�����f�u�u�;�>�3�ǫ�&����F��1������3�
�e�a�-�^��Y����]��Q��*���l�a�%�u�j�W�W���Y�Ƹ�C9��h��L���%�u�=�;��8�(���Kʹ��l_��h�E���u�d�|�0�$�}�W���Y����V
��Z�*���l�`�%�n�w�}��������l��h��L���%�u�h�}�9�8����&����R��N��ʴ�
�:�&�
�!��^����Ʈ�[��=