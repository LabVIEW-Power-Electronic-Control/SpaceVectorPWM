-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�_�&�w�8��������Z��X����_�0�!�!�w��5��=ǀ��l ��S1����g�&�f�
��(����	ӏ��F�P�����}�u�u�u�w��W���Y���	F��C����u�n�u�u�w�}�9���*����F��^ �����o�u�n�u�w�}�WϺ�ù��w2��N�����'�o�u�g�]�}�W���Y����l1��c&��U���0�0�u�h�d�f�W���Y����\��`'��=��<�!�2�'�m�}�E���Y����F�G��U�ߊu�u�u�u�;�}�W����ƿ�W9��P�����u�u�u�0�2�}�W���Y����_	��TUךU���u�u�0�u�w�}��������T��=N��U���u�<�e�u�w�3�W���&����P9��T��]���e����f�9� ���Y����F�N�����u�o�<�u�$�9��������G	��S��*����x�u�:�9�2�G��Y���F��X��U��� �u�!�
�8�4�(�������\��`'��=��1�"�!�u�~�}�W���s����V��C����=�!�6� �2�<����Ӌ��q^��sZ��E���1�
�g�&�d�3�(���J����_9��GN�����u�x�x�x�z�p�Z��T���F��Z�����x�x�x�x�z�p�Z��T���9F������;�u���f���������W��h�����%�f�u�&�w�}�W���	����l�N��U���u�4�9�u�w�}�W���Y���F��^ �����9�2�6�_�w�}�W���Y�ƭ�_��N��U���u�u�u�u�w�3�W���&����P]ǻN��U���u�u�
�-�$�<�������F���U���
�:�<�n�w�}�W���Y����l��D1�����4�u�u�u�m�4�Wϭ�����Z��R����u�:�;�:�g�f�W���Y���F��h�����!�4�<�u�w�}�MϷ�Yӕ��l
��^�U���u�u�u�u�$�<����&����RF�N��Oʼ�u�&�1�9�0�>����������Y��E��u�u�u�u�w�}��������@��h�����o�:�!�&�3�1����s���F�N�����<�
�0� �#�)����Y�ƣ�GF��S1�����#�6�:�}�f�9� ���Y��ƹF�N��N���u�0�1�6�:�2����s���K�C�X���x�x�x�x�z�����
����_F�C�X���x�x�x�x�]�}�W�������P
��N��U���!�
�:�<�l�}�Wϭ�����R��R ��U��&�1�9�2�4�W�W���������A�����u�!�
�:�>�f�W���
����_F��C
�����o�&�1�9�0�>����������Y��E��u�u�&�2�6�}�(������	F��S1�����_�u�u�<�9�1�������\��C
�����
�0�!�'�d�}�������9F������'�!�4�<�w�g��������l�N�����u�
�1�!�w�}�W���&����P9��T��]��1�"�!�u�~�W�W���������1�����u�!�
�:�>�����ۂ��9��s:��Dʱ�"�!�u�|�]�}�W�������Z��U��U���!�
�:�<��8��������d/��C����!�u�|�_�2�4�}���Y���K�C�X���x�x�x��$�<�������K�C�X���x�x�_�u�w��5��=ǀ��l��Q��*ۊ� �9�1�%�d��W�������V��Z(��M���a�
�
�%�1�9�(ށ�����@��d��Uʥ�'�u�4�u�]�}�W���Y����F�N��U���u�u�u�k�6�1�[���Y�����\��U���u�u�u�u�w�`�W�������F�N�����<�
�
�#�;�9�W���Y����l��[�����u�u�u�
�/�.�������F�S����4�4�_�u�w�}�W�������l��[��U���u�k�7�!�6�4�[���Y�����O�����4�4�u�u�w�`�W�������9F�N��U���-�&�'�&�;��������A9��V��Y���u�u�u�8�6�4�(�������W��N��U���1�!�_�u�w�f�}���Y���K�C�X���x�x�x��$�:����Y���K�C�X���x�x�_�u�w�>����Y���P
��=N��U���>�;�u�i�w�8�}���Y����R
��R��R��_�u�u�
�3�)�W��Yۂ��9��s:��Dʱ�"�!�u�u�i�z�P��������1�����u�u�<�e� ��?������\F��
P��-���u�:�u�1�9����D����Z��`'��=��1�"�!�u�w�c�P���P�Ʃ�@��^ �����n�u�u�7�#�<����D����l�N�����4�u�h�}�>�l� ���1����\��XN�H���e�|�"�0�w�u��������F�S��*����x�u�:�9�2�G��YԾ�F��EN�����7�3�u�u�w�4�F���=�����Y��E��u� �|�|�2�.�W���H����]ǻN�����u�u�i�u��9���s���K�C�X���x�x�x�x�z���������AF�C�X���x�x�x�x�]�}�W���������N�����u�u�u�u�>�}��������R��T��H��r�!�0�_�w�}�W���Y�ƥ���
N��Rʡ�0�_�u�u�w�}�W���Y�ƨ�]V��B�I���<�e�_�u�w�}�W���Y���W��h��D��u�<�d�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��d�����'�=�!�6�"�8�}