-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��LӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ��`�a�c���(���
����GF�N�����9�u�u����;���:���F��h��U���������}���Y����G��T��;ʆ�����]�}�W�������	F��cN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�%�<���6����g"��x)��N���u�<�
�0��1����Y�ƅ�5��h"��<������}�f�9� ���Y����F�^ �����4�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���)����W9��N��U���
���
��	�%���Hӂ��]��G�U���<�
�0�
�2�<�G��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����E�����u�u� �u���8���&����|4�_�����:�e�n�u�w�<�(�������\��b:��!�����
����_������\F��d��Uʴ�
�0� �;�e�g�8���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƭ�l��B��F��������4���:����U��S�����|�_�u�u�'�/����&����|3��d:��9�������w�n�W������]ǻN�����!�'�
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W�������\��yN��1�����|�_�9�f�}������P��RN�����:�u��l�f�e��������@FǻN�����4�!�4�
�8�.�(�������	F��s1��2���o�u�d�n�w�}��������R��X ��*���<�
�u�u���8���Y���A��N�����!�;�u�%���ށ�
����	F��s1��2������u�f�}�������	[�^�E��e�e�e�d�l�}�WϽ�����GF��h=�����3�8�d�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��UךU���:�&�4�!�6��#���J����lT�=��*����
����u�CϺ�����O�
N��E��e�e�e�e�g��}���Y����G����&���!�
�&�
�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�N���u�6�;�!�9�}����&����U��N�&���������W��Y����G	�N�U��e�e�e�e�f�m�G��Y����\��V ������&�c�3�:�h�Mύ�=����z%��r-��'���a�1�"�!�w�t�M���I����V��^�E���_�u�u�:�$�<�Ͽ�&����GQ��D��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��[���F��Y�����%��
�!��.�(���Y����)��t1��6���u�d�u�:�9�2�G���D����V��_�E��e�n�u�u�4�3����Y����g9��1����o������!���6���F��@ ��U���o�u�e�e�g�l�G��I���9F������!�4�
��$�l�(���&����`2��{!��6�����u�d�w�2����I����D��^�E��e�e�e�n�w�}��������R��c1��Dۊ�&�
�e�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��UךU���:�&�4�!�6��#���H����^9��T��!�����
����_������\F��T��W��d�e�e�e�g�m�U�ԜY�Ư�]��Y�����
�!�f�3�:�l�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��n�u�u�6�9�)����	����@��h��*��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I���9F������!�4�
��$�l�(���&���5��h"��<������}�c�9� ���Y���F�^�E��e�e�e�w�]�}�W���
������T�����f�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�u�W�W�������]��G1�����9�d�d�o���;���:����g)��^�����:�e�u�h�u��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�l�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�F���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�F��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��H����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������wF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����W��L�U���6�;�!�;�w�-��������9��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��_�N���u�6�;�!�9�}��������EW��T��!�����
����_�������V�S��E��u�u�6�;�#�3�W�������l
��h^��U���
���
��	�%���Y����G	�N�U��w�_�u�u�8�.��������]��[�*ٓ�o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��d�d�n�u�w�>�����ƭ�l��D�����f�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��d�e�e�w�]�}�W���
������T�����f�
��o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�d�d�g�f�W�������R��V�����
�#�g��f�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��L�U���6�;�!�;�w�-�������� 9��N��1��������}�A�������V�S��E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-��������9��N�&���������W��Y����G	�N�U��e�e�d�e�f��}���Y����G�������!�9�d�
�a�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��L�U���6�;�!�;�w�-��������9��N��1��������}�F�������V�S��E��e�e�e�d�u�W�W�������]��G1�����9�d�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����W�=N��U���&�4�!�4��2�����ԓ�\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lV�=��*����
����u�GϺ�����O�
N��E��e�e�e�w�]�}�W���
������T�����`�
�u�u���8���&����|4�]�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��u�u�6�;�#�3�W�������l
��1�U����
�����#���Q����\��XN�U��w�e�e�e�f�m�G��Y����\��V �����:�&�
�#�e��G��*����|!��h8��!���}�d�1�"�#�}�^��Y����W��^�E��u�u�6�;�#�3�W�������l
��1�U����
�����#���Q����\��XN�U��w�e�e�e�f�l�G��Y����\��V �����:�&�
�#�e�l�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�W�ߊu�u�:�&�6�)��������_��h]��3���u��
����2���+������Y��E���h�w�d�d�f�l�F��H����]ǻN�����4�!�4�
�8�.�(���A���5��h"��<������}�`�9� ���Y���F�^�E��e�e�e�e�g�f�W�������R��V�����
�#�g���g�$���5����l0��c!��]��1�"�!�u�~�g�W��H����W��L�U���6�;�!�;�w�-��������9��T��!�����
����_������\F��T��W��e�e�d�e�f�f�W�������R��V�����
�#�g���g�$���5����l0��c!��]��1�"�!�u�~�g�W��H����W��L�U���6�;�!�;�w�-��������9��T��!�����
����_������\F��T��W��e�e�d�d�f�f�W�������R��V�����
�#�
�`�m��3���>����v%��eN��U���;�:�e�u�j��F��H��ƹF��X �����4�
�:�&��+�(���Y����)��t1��6���u�`�1�"�#�}�^��Y����V��d��Uʶ�;�!�;�u�'�>��������  ��q(��3����u�u����>���<����N��
�����e�u�h�w�f�l�F��H����W��_�D��d�d�d�d�f�l�F��H����W��_�N���u�6�;�!�9�}��������EU��_��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��_�E���_�u�u�:�$�<�Ͽ�&����G9��\��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[��D��������4���Y����\��XN�U��w�e�e�e�f�f�W�������R��V�����
�#�g�f�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����W��d��Uʶ�;�!�;�u�'�>��������u#��N��1��������}�F�������V�S��D��d�d�d�d�u�W�W�������]��G1�����9�d�
�m�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��d��Uʶ�;�!�;�u�'�>��������u ��q(��U���
���
��	�%���Jӂ��]��G��H���d�d�d�d�f�l�F��H����W�=N��U���&�4�!�4��2�����ғ�\��c*��:���
�����n��������\�^�E��e�e�e�e�g�m�G��I��ƹF��X �����4�
�:�&��+�E���@����g"��x)��*�����}�d�3�*����P���W��_�E��d�n�u�u�4�3����Y����\��h��G��u�u��
���(���-���W��X����u�h�w�e�g�m�F��H��ƹF��X �����4�
�:�&��+�E���A����g"��x)��*�����}�d�3�*����P���W��_�E��e�n�u�u�4�3����Y����\��h��G��u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�d�w�_�w�}��������C9��Y����
���u�w�	�(���0����p2��F�U���;�:�e�u�j��F��H����W��_�W�ߊu�u�:�&�6�)��������_��h\�E���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����]ǻN�����4�!�4�
�8�.�(���M�ъ�u ��N��1��������}�E�������V�S��E��d�d�d�d�f�l�F��H����l�N�����;�u�%�6�9�)���&����V�=��*����
����u�DϺ�����O�
N��E��e�e�e�e�g�m�G��I���9F������!�4�
�:�$�����K����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��H����D��N�����!�;�u�%�4�3����J����\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����F��d:��9�������w�e��������\�^�E��e�w�_�u�w�2����Ӈ��P	��C1��F���o������!���6�����Y��E���h�w�e�w�]�}�W���
������T�����f�c�o����0���/����aF�
�����e�u�h�w�f��}���Y����G�������!�9�f�b�m��3���>����v%��eN��U���;�:�e�u�j��F���s���P	��C��U���6�;�!�9�e��W���-����t/��a+��:���g�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�f�W�������R��V�����
�#�
�u�w�	�(���0����p2��F����!�u�|�o�w�m�F��Y����\��V �����:�&�
�#��}�W���&����p9��t:��U��1�"�!�u�~�g�W��I��ƹF��X �����4�
�:�&��+�(���Y����)��t1��6���u�g�1�"�#�}�^��Y����]ǻN�����4�!�4�
�8�.�(���&����`2��{!��6�����u�g�3�*����P���V��UךU���:�&�4�!�6�����&����lU��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����W��^�N���u�6�;�!�9�}��������EU��X��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��_�D���_�u�u�:�$�<�Ͽ�&����G9��\��@��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�D��d�n�u�u�4�3����Y����\��h��G��u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��Y����
�c�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�d�d�e�l�}�WϽ�����GF��h�����#�g�f�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�d�e�f��}���Y����G�������!�9�g�f�m��3���>����v%��eN��U���;�:�e�u�j��F��Y����\��V �����:�&�
�#��}�W���&����p9��t:��U��1�"�!�u�~�g�W��I��ƹF��X �����4�
�:�&��+�E���Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��H����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�g�w�2����I����D��^�E��e�e�e�e�g�m�L���YӅ��@��CN��*���&�
�#�g�`��1���Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���W��_�D��d�d�d�d�f�l�F��H����l�N�����;�u�%�6�9�)���&����V��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��N�&���������W������\F��T��W��n�u�u�6�9�)����	����@��A]��E��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[�*����o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��d�e�d�d�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�f��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�l�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s�����Y������3�8�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��UךU���!�'�7�!�w�.�(�������\��C���ߊu�u�!�'�5�)�W���&����W��������3�8�o�$�:����
�Ģ�]�=N��U���;�9�4�
�>�����*����9��Z1�Oʆ�����]�}�W�������C9��P1����u�u����f�W���
����_F��G1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������z0��B��Gۊ�0�
�b�c�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������C9��P1������&�b�3�:�k�Mύ�=����z%��N�����4�u�%�&�0�?���Y�Ǝ�|*��yUךU���<�;�9�2�'�;�(��&���5��h"��<������}�f�9� ���Y����F�D������-��,�"��Fׁ�����W�=��*����
����u�FϺ�����O��N�����4�u�&�0��8�(��O����g"��x)��*�����}�u�8�3���B�����Y�����<�
�&�$���ׁ�
����	F��s1��2���_�u�u�<�9�1��������W9��T��:����n�u�u�$�:��������l ��Y�����u��
����2���+������Y��E��u�u�&�2�6�}����J����lU��N�&���������W��Y����G	�UךU���<�;�9�!�'�j����Nʹ��\��c*��:���
�����}�������9F������!�%�b�'�0�n�@���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��(�����m�
�g�o���;���:����g)��_����!�u�|�_�w�}����Ӡ��A��Y�U����
�����#���Q����\��XN�N���u�&�2�4�w��9���:���� _��G\��U���
���
��	�%���Y����G	�UךU���<�;�9����9�������
T�=��*����
����u�W������]ǻN�����9�<�8�
�"�i�F���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����'�2�f�l�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������@��h_�� ��`�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������lW��R	��M��o������!���6�����Y��E��u�u�&�2�6�}����A����_��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�n�(���&����\��c*��:���
�����}�������9F������!�%�d�b�1��Oց�H����g"��x)��*�����}�b�3�*����P���F��P ��U���
�d�
�0��e�N��*����|!��h8��!���}�b�1�"�#�}�^�ԜY�ƿ�T�������l�3�
�l��n�Mύ�=����z%��r-��'���b�1�"�!�w�t�}���Y����R
��h8��G���'�2�f�g�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����B��h��C���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϯ�&¹��T9��W��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�l�C�������F��d:��9�������w�m��������l�N�����u�
�
�d�1��Gց�K����g"��x)��*�����}�u�8�3���B�����Y�����<�
�0�
�o�m�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�d�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��Gӊ�0�
�m�`�m��3���>����v%��eN��Bʱ�"�!�u�|�]�}�W�������V
��Z�*���b�l�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��_�����m�e�o����0���/����aF�
�����e�n�u�u�$�:��������CU��Q��@ۊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����9��P1�@���u��
����2���+����W	��C��\�ߊu�u�<�;�;�4��������9��T��!�����
����_�������V�=N��U���;�9�<�8�e�/���O����`2��{!��6�����u�e�3�*����P���F��P ��U���
�l�3�
�g��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��@ӊ�0�
�m�l�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�d�<�
�"�d�F���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����g�4�9�:�2��(�������Q��N��1��������}�GϺ�����O��N�����4�u�4�2�f�<��������ZW��B1�F���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1�%���¹��_9��R��*���'�2�f�m�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������R��1�����'�&�g�<��(�N���	����`2��{!��6�����u�e�3�*����P���F��P ��U���2�d�4�9�-�/����¹��T9��V��U���
���
��	�%���Y����G	�UךU���<�;�9�%�f�m�ށ�����9��T��!�����
����_�������V�=N��U���;�9�%�d�g�4�(���&����\��c*��:���
�����}�������9F������%��9�
��(�F��&���5��h"��<������}�d�9� ���Y����F�D�����
�4�g�a�%�:�D��Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����<�
�&�$���ց�
����	F��s1��2���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������lW��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������9��E��F��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������G9��P1�D���u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&���� ^��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�o�(���&����\��c*��:���
�����}�������9F�������;�0�
�;�����K����F9��X��F��������4���Y����\��XN�N���u�&�2�4�w�<��������]��1�����f�g�u�u���8���&����|4�N�����u�|�_�u�w�4����+����9��[1�����g�<�3�
�b�o����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��<�����4�9�/�'�$�o��������F��d:��9�������w�m��������l�N�����u�0�0�0��3����&����l��N��1��������}�GϺ�����O��N�����4�u�0�0�2���������
U��N��1��������}�GϺ�����O��N�����4�u�-�
�2�0�(��&����lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�%�(�������9��E��F��u�u��
���(���-���Q��X����n�u�u�&�0�<�W����ԓ�9��h\�G���u�u��
���(���-���U��X����n�u�u�&�0�<�W����ԓ�9��P1�A���u��
����2���+������Y��E��u�u�&�2�6�}��������B9��h��E���8�l�o����0���s���@��V�����2�7�1�d�`�g�5���<����F�D�����8�
�f�
�2��N��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��#���
�e�3�
�f�n����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N��#���
�e�'�2�d�k�W���-����t/��a+��:���g�u�:�;�8�m�L���Yӕ��]��X�����
�
� �g�a��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��X�����
�
�0�
�n�k�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��S�����g�3�
�g�n�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Y
�����
�
�0�
�n�l�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��S�����g�;�!�3��o�F���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����3�:�
�
�8�����@���5��h"��<������}�w�2����I��ƹF��^	��ʥ��9�
�d�1��D���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʥ��9�
�d�%�:�D��Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����<�
�&�$����������F��d:��9����_�u�u�>�3�Ͽ�&����Q��Y�Oʗ����_�w�}����ӏ��CU��B1�E݊�g�o�����4���:����V��X����n�u�u�&�0�<�W���	����T9��V��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�e�(���K����CT�=��*����
����u�W������]ǻN�����9�!�%�m��8�(��J����g"��x)��*�����}�u�8�3���B�����Y�����!�%�e�3��i�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�`�
�0��m�G��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����g�3�
�a�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R�����
�0�
�e�`�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��A���
�a�`�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���
�e�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����Z��D��&���!�g�3�8�f�}�W���&����p]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9� ��.�4���&����P��R1�M���
�c�`�%�w�}�#���6����e#��x<��Gʱ�"�!�u�|�]�}�W�������q9��h-�����'�6� �0�f�e����M����	F��s1��2������u�e�9� ���Y����F�D�����<�;�<�
��8�(��I����g"��x)��*�����}�u�8�3���B�����Y�����9�
�e�'�0�i�C���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����
�0�
�e�f�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��Z�����b�d�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��1����`�u�u����>���<����N��
�����e�n�u�u�$�:��������9��P1�C���u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���N����lR��N�&���������W������\F��d��Uʦ�2�4�u�8��i�(���&����\��c*��:���
�����}�������9F�������;�0�
�;�����J����Q��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�6�:�E�������@9��E��A��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1�%���¹��_9��R��*���g�m�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�`�'�2�c�e�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��V ��D���9�/�'�&�c�;�(��H����	F��s1��2������u�g�9� ���Y����F�D�����4�2�d�4�;�'����M����lR��N�&���������W������\F��d��Uʦ�2�4�u�<�9�4�(݁�����
U�=��*����
����u�W������]ǻN�����9�%��9��o����M����	F��s1��2������u�d�}�������9F������$�<�
�
�2��F��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����g�3�
�m�d�-�W���-����t/��a+��:���g�u�:�;�8�m�L���Yӕ��]��C��D���'�2�a�e�w�}�#���6����e#��x<��G���:�;�:�e�l�}�Wϭ�����G��[�����a�d�u�u���8���&����|4�N�����u�|�_�u�w�4��������R��R	��D��o������!���6�����Y��E��u�u�&�2�6�}����LŹ��T9��Z��U���
���
��	�%���Y����G	�UךU���<�;�9�%��.����&����W��T��!�����
����_�������V�=N��U���;�9�%��$�1�(ہ����� R�=��*����
����u�W������]ǻN�����9�!�%�d�`�/���M����`2��{!��6�����u�e�3�*����P���F��P ��U���4�g�&�d��(�D��&���5��h"��<������}�f�9� ���Y����F�D�����
�4�g�&�f�����H���5��h"��<������}�f�9� ���Y����F�D�����%�&�2�6�2��#���H����^9��T��!�����n�u�w�.����Y����Z��S
��A���u����l�}�Wϭ�����C9��[\��C���
�g�l�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��[\��C���2�a�`�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƥ�l��t��*��� �!�'�
�`��(���J����CU�=��*����
����u�FϺ�����O��N�����4�u��6��<��������A�� _��*���
�d�m�o���;���:����g)��]����!�u�|�_�w�}����Ӈ��@��T��*���&�d�
�&��n�Mύ�=����z%��N�����4�u�%�&�0�?���H����|)��v �U���&�2�4�u��>�(�������F��E��BҊ�
� �f�e��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��{1��*���0��'�6�"�8�F���H����lR��N�&���������W��Y����G	�UךU���<�;�9�<��)�4���&����P��R1�@���3�
�a�b�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��6���
�!� �!�%��Oځ�&����W��T��!�����
����_������\F��d��Uʦ�2�4�u�0�o�;�(��L����	F��s1��2������u�g�9� ���Y����F�D�����0�m�'�2�c�j�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��{1��*���
�:�%�d�a�;�(��O����	F��s1��2������u�f�9� ���Y����F�D�����%�&�2�6�2��#���Hƹ��^9��T��!�����n�u�w�.����Y����Z��S
��B���u����l�}�Wϭ�����R��[�����:�%�g�a�e�8�G�������V��N�&���������W��Y����G	�UךU���<�;�9�0�>�>��������9��T��!�����
����_�������V�=N��U���;�9�4�'�;���������R��h��*ي� �f�g�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��3����:�
�e���(߁�&����U��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%���������C9��1�����d�3�
�c�g�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�e�i�E���H�Փ�F9��X��F��������4���Y����W	��C��\�ߊu�u�<�;�;�<����&����	��h\�*؊�
�
�
� �d�j�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��������!�%��Dف�&¹��T9��N�&���������W��Y����G	�UךU���<�;�9�6���2���+����lT��h��*���
�`�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����_��X�����g�a�g�0�f�k����K���5��h"��<������}�f�9� ���Y����F�D�����9�����)����JŹ��9��P1�B��������4���Y����W	��C��\�ߊu�u�<�;�;�>�(���<����G��h\�*���
�0�
�m�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����R��[�����:�%�g�a�e�8�G�������
_�=��*����
����u�FϺ�����O��N�����4�u��9��2�(���	����V��^��U���
���
��	�%���Y����G	�UךU���<�;�9�1�6�.��������l��N��1��������}�A�������V�=N��U���;�9�<�0�����@����	F��s1��2������u�a�}�������9F������0�%�!�%��;�(��&���5��h"��<������}�g�9� ���Y����F�D�����8�
�
� �d�h����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N�����3�
�a�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������^�����
�4�!�3��d�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
� �f�l�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�*���a�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��A���%�u�u����>���<����N��
�����e�n�u�u�$�:����&����T��h��F���%�u�u����>���<����N��
�����e�n�u�u�$�:��������lW��B1�B���u�u��
���(���-���U��X����n�u�u�&�0�<�W���&����e9��Q��Aي�a�o�����4���:����W��S�����|�_�u�u�>�3�Ϫ�	����U��]��D��������4���Y����W	��C��\�ߊu�u�<�;�;�)���M����P��G_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�:��@���&����CU�=��*����
����u�EϺ�����O��N�����4�u�
�0�"�)�@���&����CW�=��*����
����u�DϺ�����O��N�����4�u�4�
�����@����	F��s1��2������u�b�}�������9F������!�%�d�g�1��Dށ�H����g"��x)��*�����}�g�3�*����P���F��P ��U���d�3�
�l��o�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��b/��<���d�3�
�e��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���`�d�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��@���%�u�u����>���<����N��
�����e�n�u�u�$�:��������lW��B1�F���u�u��
���(���-���W��X����n�u�u�&�0�<�W���&����U��[��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.�(���&¹��@��B1�D���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&�ӓ�F9�� 1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��l�(���L�ד�F��d:��9�������w�l�W������]ǻN�����9�!�%�a��(�B���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʡ�%�a�
� �b�n����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N����
� �`�`�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h_�*���`�b�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ� 9��h[�*��o������!���6���F��@ ��U���_�u�u�<�9�1����L����lP��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�#�-�Aف�����F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_�������V�=N��U���;�9�!�%�f�e����HĹ��\��c*��:���
�����}�������9F������!�%�`�
�"�k�N���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����d�l�3�
�b��F��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��@ߊ� �c�`�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������l	��h��C���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����l ��X�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���H����P��G_��U���
���
��	�%���Jӂ��]��G�U���&�2�4�u�:��E݁�����l��N��1��������}�B�������V�=N��U���;�9�%��$�1�(݁�����l��N��1��������}�B�������V�=N��U���;�9�!�%�b����J����	F��s1��2������u�g�9� ���Y����F�D�����8�
�c�3��e�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����`�3�
�e��l�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������l ��]�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	�֓�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�F�������9��T��!�����
����_�������V�=N��U���;�9�<�8�f�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�a�
� �b�l����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����F���6�&�
�4�#�;�(��&���5��h"��<������}�f�9� ���Y����F�D�����-�
�
�
�"�i�@���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����`�
� �b�b�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��C��D���3�
�b�
�c�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������1�����m�
�g�o���;���:����g)��_����!�u�|�_�w�}����Ӗ��9��Q��L݊�g�o�����4���:����W��S�����|�_�u�u�>�3�Ϫ�	����l ��_�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�-�ށ�&����l �� W�����u��
����2���+������Y��E��u�u�&�2�6�}����I����T��G_��U���
���
��	�%���Jӂ��]��G�U���&�2�4�u�:��E���&����CT�=��*����
����u�DϺ�����O��N�����4�u��d�1��D؁�H����g"��x)��*�����}�u�8�3���B�����Y�����
� �m�d�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������9��hV�*��o������!���6�����Y��E��u�u�&�2�6�}����M����P��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�'�!����H����	F��s1��2������u�g�9� ���Y����F�D�����:�g�d�6�$����J����	F��s1��2������u�d�}�������9F������!�%�c�
�"�e�N���Y�Ɵ�w9��p'��#����u�`�u�8�3���B�����Y��'���0�
�
�
�"�e�D���Y�Ɵ�w9��p'��#����u�`�u�8�3���B�����Y�����d�3�
�m��o�Mύ�=����z%��r-��'���f�1�"�!�w�t�}���Y����R
��E1����`�<�
� �o�n����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��<�����4�9�:�0�����L����	F��s1��2������u�g�9� ���Y����F�D�����4�2�d�4�;�2����&����Q��N�&���������W������\F��d��Uʦ�2�4�u�8��j����K¹��\��c*��:���
�����}�������9F�������;�0�
�;�����&����l_��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�6�:�F�������\��h��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����]	��Q��@݊�g�o�����4���:����V��X����n�u�u�&�0�<�W���&�ޓ�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����A����
P��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)��������
9��T��!�����
����_�������V�=N��U���;�9�:�
�8�9�F؁�H����
V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9��9�8�(���&����lT��B1�@���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l ��Y�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�-�F���¹��l_��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��o�(������� 9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�F���&����CU�=��*����
����u�W������]ǻN�����9�!�%�d�d�;�(��N����	F��s1��2������u�g�9� ���Y����F�D�����8�
� �d�e��D��*����|!��h8��!���}�g�1�"�#�}�^�ԜY�ƿ�T�������!�c�3�
�g�e����Y����)��t1��6���u�`�u�:�9�2�G��Y����Z��[N�����d�3�
�e�e�-�W���-����t/��a+��:���`�u�:�;�8�m�L���Yӕ��]��C�����
�e�`�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����G��1��*��e�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����^��B1�@ߊ�f�o�����4���:����W��S�����|�_�u�u�>�3�ϳ�����F9��V��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.�(���&����l ��^�*��o������!���6���F��@ ��U���_�u�u�<�9�1����A����V��h�Oʆ�������8���L�ƨ�D��^����u�<�;�9�#�-�N���&����l��N��1��������}�B�������V�=N��U���;�9�!�%�f����N¹��\��c*��:���
�����n��������l�N�����u�8�
�e�1��F���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʡ�%�d�
� �f�l�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
� �d�b��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���d�l�
�d�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������lT��B1�Eۊ�f�o�����4���:����T��S�����|�_�u�u�>�3�Ϫ�	����U��]�����u��
����2���+������Y��E��u�u�&�2�6�}����A����G9��h_�D���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&�ԓ�F9��^��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������S��N�&���������W������\F��d��Uʦ�2�4�u�8��k����H�ӓ�F��d:��9�������w�l�W������]ǻN�����9�!�%�f��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�d�
� �f�j�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����� �d�m�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��]�� ��m�
�f�o���;���:����g)��[�����:�e�n�u�w�.����Y����^��B1�Lފ�d�o�����4���:����S��S�����|�_�u�u�>�3�Ϫ�	����U��W�����u��
����2���+������Y��E��u�u�&�2�6�}�(�������l ��\�*��o������!���6��� F��@ ��U���_�u�u�<�9�1����Hƹ��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Fׁ�����9��T��!�����
����_�������V�=N��U���;�9�%��;��(���H����CU�=��*����
����u�DϺ�����O��N�����4�u�8�
�d�;�(��I����	F��s1��2������u�g�9� ���Y����F�D�����
� �d�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��^1�����g�a�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӗ��U��[�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�,�(�������l ��\�*��o������!���6�����Y��E��u�u�&�2�6�}����I����T��h�Oʆ�������8���K�ƨ�D��^����u�<�;�9�'��݁�&����S��G\��U���
���
��	�%���Jӂ��]��G�U���&�2�4�u�:��(���H����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'����N����\��c*��:���
�����}�������9F������&�9�!�%��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�c�
� �f�o�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�d�3�
�e�n����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���b�3�
�g�c�-�W���-����t/��a+��:���g�u�:�;�8�m�L���Yӕ��]��D�����f�3�
�g�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����
� �d�e��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�g�l�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��[1�����3�
�f�b�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������hX�� ��m�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����G�� 1��*��g�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������9��h_�M���u�u��
���(���-���U��X����n�u�u�&�0�<�W���&����9��h_�L���u�u��
���(���-���U��X����n�u�u�&�0�<�W���&�Г�F9��X��F��������4���Y����\��XN�N���u�&�2�4�w�0�D�������T��Q��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	¹��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'�.�(���H����CT�=��*����
����u�FϺ�����O��N�����4�u�:�g�1��D���	����`2��{!��6�����u�d�w�2����I��ƹF��^	��ʡ�%�m�
� �f�e�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��ۊ�4�!�3�
�d�d����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N����
� �d�e��l�Mύ�=����z%��r-��'���f�1�"�!�w�t�}���Y����R
��Z��C���
�a�a�%�w�}�#���6����e#��x<��@���:�;�:�e�l�}�Wϭ�����_"��B1�Dڊ�d�o�����4���:����V��X����n�u�u�&�0�<�W���&���� _��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'����Hǹ��\��c*��:���
�����}�������9F������!�%�d�m�1��C���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�b�3�
�c�m����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����D���
�a�a�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������\��T��*���d�c�
�d�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������^��1��*��g�%�u�u���8���&����|4�]�����:�e�n�u�w�.����Y����VT��h_�� ��`�
�g�o���;���:����g)��[����!�u�|�_�w�}����Ӕ��l ��Z�*��o������!���6��� F��@ ��U���_�u�u�<�9�1��������9��Q��A���%�u�u����>���<����N��S�����|�_�u�u�>�3�ό�����R
��X ��*���d�c�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�d�<�3��i�C���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����d�4�9�:�2��(���H����CT�=��*����
����u�W������]ǻN�����9�!�%�f��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʇ�;�0�
�9��8��������9��T��!�����
����_�������V�=N��U���;�9��;�2���������9��h_�M���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Kʹ��G9��h_�E���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����J¹��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����A����S��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����R��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�:��2���&����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9��3�ށ�����V��B1�MҊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����9��h_�M���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1���@����F9��Z��G��������4���Y����\��XN�N���u�&�2�4�w��E݁�&����V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)��������R��N�&���������W������\F��d��Uʦ�2�4�u�0��0�Bہ�����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�(���H����CT�=��*����
����u�W������]ǻN�����9�6�'�,�f�3��������
T��N�&���������W������\F��d��Uʦ�2�4�u�4�0�o��������9��C1�����`�m�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lW��h��D��
�f�o����0���/����aF�
�����e�n�u�u�$�:��������VW��h�� ��e�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����VW��[�����g�8�-�<�1��A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���g�
�
� �f�o�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*���<�;�f�3��k�O���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����b�3�
�c�e�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��G1��؊�
� �d�a��o�Mύ�=����z%��r-��'���b�1�"�!�w�t�}���Y����R
��R����
� �d�`��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�c�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��Fߊ� �d�b�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��F���
�c�f�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����@��C��C���
�c�e�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����G��\�����c�d�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ�� W��S�����
� �d�l��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��GY�� ��l�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����_T��1��*��m�%�u�u���8���&����|4�Y�����:�e�n�u�w�.����Y����J9��^_�� ��e�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����G��^����� �d�g�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������9��C1��*���d�f�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�d�;�!�>����M����\��c*��:���
�����}�������9F������7�8�'�0�e��F���&����l��N��1��������}�GϺ�����O��N�����4�u�4�2�f�<��������^��^_�� ��`�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����VW��[�����g�<�
�`�1��@���	����`2��{!��6�����u�e�3�*����P���F��P ��U���0�0�
�;�$�l����N�ޓ� F��d:��9�������w�m��������l�N�����u�0�
�8�c����NŹ��\��c*��:���
�����}�������9F������;�"�<�;�>��(���H����CU�=��*����
����u�W������]ǻN�����9�!�%�e�1��@���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�a�
�"�l�Nׁ�K����g"��x)��*�����}�u�8�3���B�����Y�����c�
� �d�`��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����f�3�
�b�d�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R�����0�:�
�
�"�l�Fց�J����g"��x)��*�����}�u�8�3���B�����Y�����!�1�/�'�$�l��������V��N�&���������W������\F��d��Uʦ�2�4�u�0�2�8�(�������]	��^_�� ��d�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����A��^_�� ��g�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����W��B1�G݊�g�o�����4���:����V��X����n�u�u�&�0�<�W�������\��h^��D���
�b�d�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������A��P�D���8�'�4�
�f�;�(��A����	F��s1��2������u�g�9� ���Y����F�D�����<�;�4�&�0��(���H����CU�=��*����
����u�W������]ǻN�����9�7�8�'�2�o�(�������R��N�&���������W������\F��d��Uʦ�2�4�u�;�2�;����&����S��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�:�2�;����&����U��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�0������ד�\��B1�C؊�g�o�����4���:����V��X����n�u�u�&�0�<�W���H¹��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�5�0��������U��[�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����_��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�%��1�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�0��0�F�������T��Q��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����S��B1�Eڊ�f�o�����4���:����W��S�����|�_�u�u�>�3�ϼ�����9��h_�A���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l ��W�*��o������!���6�����Y��E��u�u�&�2�6�}���&����
T��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)�������� W��N�&���������W������\F��d��Uʦ�2�4�u�
�6�o�F߁�����lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�8�(���MŹ��lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�<��������]��1��Dފ� �d�a�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��G���
�l�l�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��Q��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����R��B1�Bӊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&�Փ�F9��]��G��������4���Y����\��XN�N���u�&�2�4�w�8�(���K����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�3�1��������l ��W�*��o������!���6�����Y��E��u�u�&�2�6�}��������A	��Y�����l�d�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӂ��V��h�����
�:�
�
�"�l�N؁�K����g"��x)��*�����}�u�8�3���B�����Y�����'�0�<�3��m�E���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����`�3�
�e�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R�����;�&�e�<�1��N���	����`2��{!��6�����u�e�3�*����P���F��P ��U���0�2�d�d�3�0����&����lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�:�(�������F9��]��F��������4���Y����\��XN�N���u�&�2�4�w�/����H�ד�l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}��������U��\�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�2��������lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�:�(�������\��B1�Aۊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���L����V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�%�8����&����lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�D݁����� 9��T��!�����
����_�������V�=N��U���;�9�%��;��(���K����CU�=��*����
����u�DϺ�����O��N�����4�u�0�
�:�d�(�������l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}��������U��Y�����u��
����2���+������Y��E��u�u�&�2�6�}��������lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����N����V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:�k����H�ד�F��d:��9�������w�m��������l�N�����u�0�
�8�e����IĹ��\��c*��:���
�����}�������9F������%��9�
��(�(���K����CU�=��*����
����u�DϺ�����O��N�����4�u�0�
�:�o�(���K����CU�=��*����
����u�DϺ�����O��N�����4�u�
�4�e�o�(���J����CT�=��*����
����u�CϺ�����O��N�����4�u�8�
�d����Lǹ��\��c*��:���
�����}�������9F������!�%�d�l�1��F���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
� �g�`��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��^1��*���g�b�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƽ�Z��B1�A݊�f�o�����4���:����V��X����n�u�u�&�0�<�W�������]9��Q��D���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϯ�/����_��B1�FҊ�a�o�����4���:����T��S�����|�_�u�u�>�3�Ϫ�	����U��V�����u��
����2���+������Y��E��u�u�&�2�6�}��������lT��B1�Lӊ�f�o�����4���:����V��X����n�u�u�&�0�<�W���&����U��X�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�%��.����M����l ��\�*��o������!���6�����Y��E��u�u�&�2�6�}��������lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�9�)���� ����T��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�6�/�(���K����CT�=��*����
����u�W������]ǻN�����9�1�9�!�3�'����K����T��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��2�(�������
9��T��!�����
����_�������V�=N��U���;�9�7�8�%�8�݁�����9��T��!�����
����_�������V�=N��U���;�9�!�%�`����JĹ��\��c*��:���
�����}�������9F������%�f�
�
�"�o�C܁�K����g"��x)��*�����}�u�8�3���B�����Y�����'�0�e�1�:�/����&����P��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�l�(�������l ��\�*��o������!���6�����Y��E��u�u�&�2�6�}���&����^��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�j�(���K����CT�=��*����
����u�W������]ǻN�����9�3�%�������
����V9��[��L݊�
� �g�e��o�Mύ�=����z%��r-��'���f�1�"�!�w�t�}���Y����R
��E�����
�g�3�
�d�d����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������g�
� �
�"�o�E܁�J����g"��x)��*�����}�f�3�*����P���F��P ��U���4�g�d�3��n�G���Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����d�d�3�
�d�n����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���3�
�f�b�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W������� ��h/�����
�7�:� �2�����@ʹ��U��X�����u��
����2���+������Y��E��u�u�&�2�6�}����;����G9��D�����4� �
�b�f�;�(��K����	F��s1��2������u�e�}�������9F������3�%����)�6�������e��R1�*ۊ� �g�c�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��G��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������t#��B�����0�
�'��"�1����&����l��N��1��������}�GϺ�����O��N�����4�u�:�9�/��8���>����V��E1�� ���d�3�
�f�f�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��X������!��0�#�/�8�������@9��h\�B���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����H�ԓ�F9��W��F��������4���Y����\��XN�N���u�&�2�4�w�0�(�������_��N�&���������W������\F��d��Uʦ�2�4�u�0�`�;�(��J����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�a��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʼ�8�f�
�:��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�b�
� �e�l�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�d�3�
�c�l����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���d�`�1�8�%�<�(���K����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�e�(�������l ��Z�*��o������!���6�����Y��E��u�u�&�2�6�}����I����R��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����Q��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�3�'�3��������V��h��G��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������\��C��*��
�
� �g�g��F��*����|!��h8��!���}�a�1�"�#�}�^�ԜY�ƿ�T����*���0�!�'�
�g��(���K����CT�=��*����
����u�CϺ�����O��N�����4�u�'�6�9����HŹ��\��c*��:���
�����}�������9F������;�"�0�
�"�o�E߁�J����g"��x)��*�����}�a�3�*����P���F��P ��U���6�;�d�3��h�@���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����;�g�3�
�b�d����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�� ��&���
� �g�f��n�Mύ�=����z%��r-��'���a�1�"�!�w�t�}���Y����R
��O�����!�'�
�l�����@ǹ��\��c*��:���
�����i��������l�N�����u�0��9��(�E��&���5��h"��<������}�c�9� ���Y����F�D�����0��9�
�"�o�A؁�J����g"��x)��*�����}�a�3�*����P���F��P ��U����9�
� �e�k�(��Cӵ��l*��~-��0����}�a�1� �)�W���s���@��V�����9�
� �g�n��D��*����|!��h8��!���}�f�1�"�#�}�^�ԜY�ƿ�T�� ��&���a�
�4�!�1��B���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʻ�"�0�c�3��k�@���Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����0�g�3�
�a�m����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N�����%�`�3�
�a�n����Y����)��t1��6���u�g�1�"�#�}�^�ԜY�ƿ�T����*���g�e�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G[�����c�m�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��X�� ��f�
�f�o���;���:����g)��\�����:�e�n�u�w�.����Y����_T��h��G��
�f�o����0���/����aF�N�����u�|�_�u�w�4����	����9��Q��@���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l ��X�*��o������!���6���F��@ ��U���_�u�u�<�9�1����A����lT��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�����L����U��Y�����u��
����2���+������Y��E��u�u�&�2�6�}�(���K����U��Z�����u��
����2���+������Y��E��u�u�&�2�6�}����O����P��h�Oʆ�������8���K�ƨ�D��^����u�<�;�9�#�-�Oځ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�
�����O¹��\��c*��:���
�����h��������l�N�����u�-�
���$��������_��Z��*���g�m�
�e�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������^��1��*��`�%�u�u���8���&����|4�X�����:�e�n�u�w�.����Y����K+��c�����9�<�9�
�e��(���K����CW�=��*����
����u�BϺ�����O��N�����4�u�
�
��(�E��&���5��h"��<������}�b�9� ���Y����F�D�����-�
���.�(�(�������lW��h8�� ��l�
�e�o���;���:����g)��]����!�u�|�_�w�}����Ӏ��l��{:�� ��� �!�%�,�f�j�!���&����l��N��1��������}�E�������V�=N��U���;�9�3�%�/��#�������G��N1�A���3�
�c�l�'�}�W���&����p9��t:��U���u�:�;�:�g�f�W���
����_F��e�����
�b�3�
�`�d����Y����)��t1��6���u�d�1�"�#�}�^�ԜY�ƿ�T�������!�d�3�
�`�h����Y����)��t1��6���u�g�1�"�#�}�^�ԜY�ƿ�T����*����,� �
�"�)����H�ѓ�l ��X�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������_��N�&���������W������\F��d��Uʦ�2�4�u�
��n����A�ғ�F��d:��9�������w�m��������l�N�����u�7�4�&�0��(���K����CT�=��*����
����u�W������]ǻN�����9�!�%�l��(�E��&���5��h"��<������}�f�9� ���Y����F�D�����
�4�g�`��(�E��&���5��h"��<������}�f�9� ���Y����F�D�����0�&�2�7�#�n����@�Փ� F��d:��9�������w�m��������l�N�����u�8�
�d�1��N���	����`2��{!��6�����u�e�3�*����P���F��P ��U���'�
�
� �e�l�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
� �g�g��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��_��D���
�l�f�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��R
�����
�
� �g�e��D��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��G1�����
� �g�`��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��Z�����
� �g�`��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���g�c�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƨ�_��S1�����
� �g�f��n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��V��D���
�l�`�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������A��P�*���:�2�;�<��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�g�
�0�8�:����&����l��N��1��������}�GϺ�����O��N�����4�u�8�d��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʠ�1�'�9�"�d�;�(��H����	F��s1��2������u�g�9� ���Y����F�D�����#�'�9�"�d�;�(��N����	F��s1��2������u�g�9� ���Y����F�D�����8�d�
� �d�m�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����0�<�<�
�"�o�Nف�K����g"��x)��*�����}�u�8�3���B�����Y�� ���'�9�"�f�9�)����I�ޓ�F��d:��9�������w�m��������l�N�����u�
�4�g�e�l��������R��N�&���������W��Y����G	�UךU���<�;�9�%��1�(݁�A���� V��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�%�i����I�ޓ�F��d:��9�������w�m��������l�N�����u�
�
�a�1��G���	����`2��{!��6�����u�e�3�*����P���F��P ��U���4�&�2�
��(�D��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�l�
� �d�h�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*���g�`�
� �d�h�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����2�7�!�a�1��G���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�`�3�
�g�m����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������
� �f�b��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��Y	��*���
�;�&�c�1��G���	����`2��{!��6�����u�e�3�*����P���F��P ��U���2�d�4�9�-�/��������
W��N�&���������W������\F��d��Uʦ�2�4�u�4�0�o��������9��h]�D���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����@Ź��lU��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'�i�(�������_��N�&���������W������\F��d��Uʦ�2�4�u�0�2�8�(�������U��W�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�-��������lU��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�5�0����ǹ��lU��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�N؁�����9��T��!�����
����_�������V�=N��U���;�9�1�9�#�9����&����lU��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'�n�(�������U��N�&���������W������\F��d��Uʦ�2�4�u�'�2�:�C߁�����R��1��*��g�%�u�u���8���&����|4�N�����u�|�_�u�w�4�������� 9��Z����� �f�`�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��1��*��a�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������U
��hZ�� ��b�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����U
��hZ�� ��a�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����9��h]�D���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l��Q��D���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϫ�����\��h ��*���f�m�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƽ�e��h\�*���
� �f�l��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��h8��G���g�
� �f�g��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����DҊ� �f�d�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������Y��*���8�d�e�3��o�F���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����l�
� �f�e��C��*����|!��h8��!���}�e�1�"�#�}�^�ԜY�ƿ�T�������4�0��'�4�(���A���� T��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�>�����
����A��B��D���3�
�g�e�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�*���f�`�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��1��*��`�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��h��F��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CT��h
�����;�3�
�g�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��Eۊ� �f�c�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��E���
�g�m�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�E���8�'�4�
�"�n�G߁�K����g"��x)��*�����}�u�8�3���B�����Y�����d�g�3�
�e�h����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���c�
� �f�g��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����f�3�
�f�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����
� �f�l��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�g�c�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������T������'�6� �2�l�B���&����l��N��1��������}�D�������V�=N��U���;�9�:�
�8�9�(���J����CT�=��*����
����u�W������]ǻN�����9�;�"�0�`�;�(��A����	F��s1��2������u�d�}�������9F������;�"�0�m�1��D���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʺ�
�:�1�
�"�n�C߁�K����g"��x)��*�����}�u�8�3���B�����Y�����:�1�
� �d�k�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����d�
� �f�b��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�� ��&���e�3�
�f�a�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��Y����
� �f�b��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��R�����3�
�f�f�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��@=��Dߊ� �f�l�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������d��A���
�f�d�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����]��R�*���f�d�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������V��[_�����a�l�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƣ�D5��Y�� ��g�
�f�o���;���:����g)��]����!�u�|�_�w�}����ӏ��_��X�����g�d�3�
�c�o����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N����l�3�
�a�g�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��Cڊ� �f�l�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��[�����a�d�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�Z*��C1�����:�
�
� �d�m�(��Cӵ��l*��~-��0����}�e�1� �)�W���s���@��V�����e�
� �f�`��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����3�
�`�d�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������{1��*���
�:�%�6�$����Hù��\��c*��:���
�����l��������l�N�����u�;��'�8��(�������A9��X��*���f�d�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������V
��Z�����`�a�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��1��*���e�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��Q��@���%�u�u����>���<����N��
�����e�n�u�u�$�:�����ߓ�F9��V��G��������4���Y����\��XN�N���u�&�2�4�w�8�(���O���� S��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2���������S��N�&���������W��Y����G	�UךU���<�;�9�<��8�ށ�����T��Y
�����0�g�3�
�b�j����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*�����!�g�n�;�(��L����	F��s1��2������u�d�}�������9F������!�%�d�a�1��B���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʴ�'�9�
�:��2���M�֓�lV��B1�Mڊ�d�o�����4���:����U��S�����|�_�u�u�>�3�ϭ�����9��h]�E���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l ��X�*��o������!���6�����Y��E��u�u�&�2�6�}��������l*��G1�A���0�e�3�
�b�k����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����
�:�
�:�'�o�C����֓�l ��X�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������A9��X��Eފ�
�
�
� �d�e�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����!��'��8��Gہ�&����U��Z�����u��
����2���+������Y��E��u�u�&�2�6�}��������l*��G1�A���0�d�g�3��k�O���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����9�
�b�3��j�O���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����3�
�g�
�2�g�$���5����l�N�����u�%�&�2�4�8�(���
�ԓ�@��T��!�����n�u�w�.����Y����Z��S
��E��o�����W�W���������D�����
��&�f�1�0�E��*����|!��d��Uʦ�2�4�u�%�$�:����K����	F��x"��;�ߊu�u�<�;�;�<�(���&����l5��D�����f�o�����4�ԜY�ƿ�T�������7�1�g�e�w�}�8���8��ƹF��^	��ʴ�
�<�
�&�&��(���&����F��d:��9����_�u�u�>�3�Ͽ�&����Q��_�U������n�w�}�����ƭ�l��h�����
�!�
�&��}�W���&����p]ǻN�����9�4�
�<��9�(��J����|)��v �U���&�2�4�u�%����N����	F��s1��2���_�u�u�<�9�1��������lV��E��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��n�u�u�&�0�<�W�������]9��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�>�3�Ͽ�&����A��h����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�n�u�u�$�:����	����F��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4��������G��hZ�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�.����Y����V��Y1�����u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}����Ӈ��}5��D��U���
���
��	�%���Mӂ��]��G�U���&�2�4�u�'�.��������F��u!��0���_�u�u�6�:�2��������R��Q1�����
�g�&�f�9��E��0���F��Y�����u�u�u�u��}�W���<����9F�N��U���
���u�w��2���B���F�
��E�����o����%�ԜY���F��Y_��<���u�u����f�W���Y����\��`'��=������~�W�W������9F�N��U���u�u�����0���s���F�E�����u��
���L���Y�����N�<����
�����#���Q����\��XN�N���u�u�u�1�9�}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY���F��T��;ʆ�����]�}�W���Y����\��b:��!�����
����_������\F��G�U���0�1�6�8�8�8��Զs���P	��X ��ʸ��`�a�c������&�Ԣ�lP��N�����u�0�0�<�w�W�W���Y�ƅ�\��y:��0��u�u�u�u���$���<����}2��r<�U���u�u�1�;���#���Y����t#��=N��U���u�:�!����Mϗ�-����O��N�����u�_�u�u�w�}���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF�N�����o������0���/����aF�N�����u�|�|�_�w�}��������V��=dךU���:�%�;�;�w��N��Aŀ��l��h]��D���9�
�g�d��W�W�������PF�N��U����u�u����L���Y���(��h=��2���u����l�}�W���Yӂ��9��s:��Oʜ����_�w�}�W����ԓ�z"��T��;����n�u�u�w�}����&����{F��~ ��2���_�u�u�u�w�4�C���=���/��r)��N���u�u�u�1�"��>���Y�ƅ�g#��eN����u�:�!�}�w�}�W�������	F��=��*����
����u�FϺ�����O��N��U���1�;�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���Y����\��yN��1��������}�D�������V�=N��U���u�<�a�o��}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W���Y����\��b:��!�����
����_������\F��G�U���0�1�6�8�8�8��Զs���P	��X ��ʸ��`�a�c����������]����@���_�u�u�2�8����s���F�~*��U�����n�u�w�}�Wϐ�4����t#�'��0���n�u�u�u�w�9�߁�0����	F��c+��'�ߊu�u�u�u�>�l� ���1����}2��r<�U���u�u�1� ���#���Y����t#��UךU���:�!�}�u�w�}�WϺ�����z(��c*��:���
�����k��������l�N��Uʱ�;�u�u����;���:����g)��_����!�u�|�_�w�}�W������)��=��*����
����u�CϺ�����O�d��Uʰ�1�6�8�:�2�)�}�Զ����9F���*���#�f�;�
�e�.�D݁�&�����G������l�d�m�1�m����&�Ԣ�lU��D1�*�ߊu�u�0�0�>�}����s���F�~*��K��_�u�u�u�w��(���>���Q�N��U���1�;�
���}�I��U���F�
��D�����h�u�e�W�W���Y�ƨ�F��~*��U��f�|�u�u�'�/�W���Y���F�N����u�%�6�>�]�}�W���Y����GF������_�u�u�u�w�4�G��Y����V ��[��*���u�u�u�u�3�3�W�������U9��O1����u�u�u�0�j�}��������l��=N��U���u�:�!�h�w�/�(���J�ד�O��=N��U���
�1�#�f�9��E���J����fW������;�u��l�f�e�������� T��h]����
�_�u�u�2�8�������F�N��<���k�d�_�u�w�}�W���&����vF�Y�U���u�u�1�;���#���G����9F�N��U���d����j�}�E�ԜY���F��B��<���u�k�f�|�w�}����Y����l�N��Uʶ�>�h�u�%�4�6�}���Y���A��CN��U���'�!�_�u�w�}�W���I���Z��R�����e�_�u�u�w�}���D�ƥ�l��h��*���u�u�u�u�4�}�IϹ�	���� T��T�U���u�u�1� �w�c��������9��UװU���3�e�3�0�#�n����M�ד�F��T�����!�8��`�c�k�(߁�	���� T��hX��D���u�2�;�'�4�0����Y���F��sN��U���u�u�u�u���$���<���JǻN��U���<�e����`�W��s���F�S��*����u�k�c�~�}�WϮ��ơ�CF�N��U���1�;�u�k�1��3���6����W��R	��B��_�u�u�u�w�2���Y����@��h��F���%�|�_�u�w�;�G���������Z��*��o�6�8�:�2�)����L����U9��Q����;�
�a�d�w�}��������R�=N��U���u��h�u�{�}�W���YӨ��l5��p+��K��_�u�u�u�w�4�G���=���F��d��U���u�1� �
��	�W���O��ƹF��X�����}�u�u�u�w�9����GӀ��K"��N!��*��
�0�
�b�f�W�W���Y�ƨ�F�	N�����2�
�
� �d�k����s��� ��h��*١�d�&�9�
�e�l�"���Y����\��CN��3���a�c�
�
�"�����
���� T��=N��U���0�<�u�4�w�W�W���Y�ƅ�[�BךU���u�u� �
���W���H���F�N��ۊ���u�k�d�q�W���Y����Z��`'��=��u�g�_�u�w�}�W���J����g.�	N�Y���u�u�u�1�9��>���Y���l�N��Uʱ� �
���w�c�D���Y����\��Z��]���u�u�u�1�9�}�IϷ�&����R��d�����0�d�`�f�%�:�C��U���F�
��G��u��6�
�6�8�$�������lW��h_�����d�f�_�u�w�}�W���J���Z*��C1�����!� �!�'��j�(݁�����^�N��U���1�;�u�k�>���������C9��E��F��_�u�u�u�w�2���Y����G9��E1�����e�
� �f�a��B��s���U9��Z�����d�;�
�m��h�F���Y�Ư�^��R �����`�a�c�
��(�(���&�Ѣ�lW��h]��D���u�2�;�'�4�0����Y���F��sN��U���u�u�u�u���$���<���JǻN��U���<�e����`�W��s���F�S��*����u�k�d�{�}�W���Yӂ��G9��s:��H���`�_�u�u�8�)����Q���F�
��E��u�
�4�g�e����H˹��l�N��Uʱ�;�u�k�3�'�)����K�ғ�l��h]�D�ߊu�u�u�u�8�)�J���&����lT��Q��B���%�|�_�_�]�}�W��Y����P��R �����0�}�%���.�^ϱ�Y����@��RN�����0�u�x�u�w�<�(�������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N�����
�&�u�h�6��#���H����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�&�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����0� �;�e�'�8�W�������A	��D�X�ߊu�u�%�'�#�/�(߁�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N�����!�'�
�
�%�:�K���	����@��A]��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(��Y����]	�������1�3�
�a�g�-�W���	����@��A_��\���u�=�;�_�w�}�W���Y���F�N��*��� �;�e�%�2�}�JϿ�����u	��{��*��
�
�
�
��8�(��B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�4��8����H����TF��D��U���6�&�{�x�]�}�W�������]9��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�%�%�)����&����Z�V�����
�#�g�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���Hƹ��^9��N��ʻ�!�}�-�!�8�9����M�֓�F�V�����
�#�
�|�~�}����s���F�N��U���u�u�4�
�2�(����	����[��E�����'��:�
�g��(���&Ź��T9��UךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W������G��h\�����4�&�2�u�%�>���T���F��h�� ���g�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���	����F��1�����h�4�
�:�$�����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C_�����d�|�4�1�9�)�_�������l ��Z�*��h�4�
�:�$��ށ�P���G��d��U���u�u�u�u�w�}�WϿ�&����A��h����u�9��������&����V9��E��G��_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����E�����
�'�2�4�$�:�W�������K��N�����0� �;�f�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���R��R�����%�0�u�h�6�����&����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���`�3�8�d�~�<�ϰ��Ω�Z��Y
�� ��`�
�g�h�6�����&����O�N�����u�u�u�u�w�}�W���Y����C9��C��*ي�'�2�i�u�;��3���+����^9��1��D���2�g�`�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C�����!�'�
�
�%�:�����Ƽ�\��D@��X���u�4�
�0�"�3�C�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��*��� �;�a�%�2�}�JϿ�&����G9��\��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�`�1�0�F�������\�R�����
� �f�`��o�JϿ�&����G9��1�\���!�0�u�u�w�}�W���Y���F������'�
�
�'�0�a�W���0����r4��R��G���0�e�'�2�e�j�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�%�'�!�%��(���Ӈ��Z��G�����u�x�u�u�6������ӓ�A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���4�
�0� �9�h����Y����C9��Y����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�B��������� ��]°�<�6�;�
�"�n�B߁�K����C9��Y�����e�|�|�!�2�}�W���Y���F�N��U���%�'�!�'������E�Ư�l/��r6��'���8�g�c�0�f�/���M���F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u��1�(���&����l��R	��D���&�<�;�%�8�8����T�����[�����:�%�&�'�0�n�G���
����C��T�����&�u�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��R���=�;�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�3�}�'�.��������O��_�����u�u�u�u�w�}�W���Y����Z9��E1�����
�0�
�d�w�`��������l*��G1�C���
�a�c�%�l�}�W���Y���F������}�%�6�;�#�1����H����C9��P1������&�d�
�$��D�������9F�N��U���u�u�u�u�w���������\��h��*��u�h�4�
�8�.�(���&��ƹF�N��U���u�u�;�u�1�W�W���Y���F��SN��N�ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠu�u�x�u�$�4�Ϯ�����F�=N��U���6�&�u�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��R��u�=�;�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1����|�u�=�;�w�}�W���Y���F��1����b�u�h���(�D���	��ƹF�N��U���u�u� �������J����[��b/��<���3�
�l�
�e�W�W���Y���F�N�����
�9�
�;�$�o�ށ�����W�
N�����
�9�
�;�$�o�ށ�����l��=N��U���u�u�u�u�w�<��������V��h\��D���2�f�m�u�j�����&����I��D1��ۊ� �l�l�%�l�}�W���Y���F�<�����4�9�:�0���F�������F�<�����4�9�:�0���F���&����CU��N��U���u�u�u�u�>�0�E������� F���؊� �b�d�%�l�}�W���Y���F������2�f�l�u�j�4��������l��=N��U���u�u�u�u�w�.����&���� ^��R�����
�
�
� �c�j����Jӂ��]��]����u�u�u�u�w�}�W�������T9��X��Hʼ�0�
�
� �d�d����Jӂ��]��]����u�u�u�u�w�}�W���Kù��l��h]�F��u�
�g�
�f�;�(��L����9F�N��U���u�u�u�
�6�o�N�������F������l�3�
�l��n�}���Y���F�N�����
�0�
�m�n�a�W���H����T��G]�U���u�u�u�u�w�}����¹��T9��^��Hʧ�<�<�
� �`�d���Y���F�N��U���0�
�8�g��8�(��L���@��C��L���
�d�
�f�]�}�W���Y���F�D�����d�'�2�f�b�}�Jϭ����� W��B1�L���n�u�u�u�w�}�W���Yӕ��l��Y�����m�c�i�u�2����&����W��UךU���u�u�u�u�w�}����HĹ��T9��W��Hʡ�%�d�b�3��e�(��s���F�N��U���!�%�d�a�%�:�D��Y����l0��1�����l�
�f�d�w�2����H����F�N��U���u�u�!�%�f�����N���F��G1�*���f�`�%�n�w�}�W���Y���F��Z��M���2�f�d�u�j�)���&����
U��UךU���u�u�u�u�w�}����@����lU��N�U���
�l�3�
�g��E�ԜY���F�N��Uʡ�%�b�'�2�d�j�W������l ��Y����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��ƓF�C�����;�%�:�0�$�}�Z���YӖ��P��F��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y�����Yd��U���u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���ց�
����O��_��U���u�u�u�u�w�}�%���¹��_9��R��*���0�
�l�`�k�}����H����l	��D1�����
�`�c�%�l�}�W���Y���F�<�����4�9�/�'�$�o��������F�<�����4�9�/�'�$�o����&����l��=N��U���u�u�u�u�w�<����&����T9��[��Hʶ�'�,�d�<�1��D���	��ƹF�N��U���u�u�0�0�2���������
U��S�����0�
�;�&�1��A���	��ƹF�N��U���u�u�-�
�2�0�(��&����T9��_��Hʳ�%�!�'�g�e�i�!���&����l��=N��U���u�u�u�u�w�8��������V��_�I���
�4�g�a�1��D���	������Y��G���_�u�u�u�w�}�W���Y����_T��h��*��m�i�u�
�6�o�C���&����l��=N��U���u�u�u�u�w�0�(�������
W��S�����g�3�
�f�g�-�L���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�u�u�x�w�.����	����@�CךU���'�6�&�u�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H��r�u�=�;�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�d�|�u�?�3�W���Y���F�N�����d�4�9�:�2��(���&����Z�e��ۊ�9�
�;�&�b�;�(��L����9F�N��U���u�u�u�4�0�l��������lR��R	��E��i�u�4�2�f�<��������l ��Y�*��_�u�u�u�w�}�W���Y����VT��[�����f�'�2�a�`�}�Jό�����R
��X ��*ي� �g�c�
�e�W�W���Y���F�N��'���9�
�
�0��l�N��Y����K+��c�����9�<�9�
�e��(���K����CT�N�����u�`�n�u�w�}�W���Y�����R�����'�2�a�f�w�`��������J)��h#�����,�d�b��1��A���	������Y��@���_�u�u�u�w�}�W���Y����_T��1����a�u�h�3�'�%�"���6����F
��G��D����3�
�c�n�-�_������\F��UךU���u�u�u�u�w�}�(���K����A��^�U��3�%�-� ����������J9�� 1�����c�l�%�}�d�9� ���Y���9F�N��U���u�u�u�7�#�l����M����[��O��8���,� �
� �#�-���M����F9��W��G��u�:�;�:�e�t�}���Y���F�N�����
�
�0�
�f�i�K�������f*��x��8���<�9�
�g�����@ʹ��T��S�����d�n�u�u�w�}�W���Y����Z��^��*���
�e�e�i�w�%�(���5����G9��[�����g�
�
� �e�e�(��L�ƨ�D��[�N���u�u�u�u�w�}�Wϭ�����lT��R	��E��i�u�-�
������&����Z��h_�*��� �g�l�
�e�h�W������O��N��U���u�u�u�u�#�-�F�������S��S�����a�
� �g�d��F�ԜY���F�N��Uʡ�%�d�c�'�0�i�A���DӀ��l��{:�� ��� �!�%�,�f�i�!���&����l��]�����:�`�|�_�w�}�W���Y���F��G1�B���2�a�c�u�j�;����,����F��B�����d�a��3��k�N���Q����\��XN�\�ߊu�u�u�u�w�}�W�������
9��P1�B���h�3�%�-��	�8���4����C
��\��#���
�c�l�%��i��������]ǻN��U���u�u�u�u�:��B݁�����_�
N����g�3�
�m�d�-�L���Y���F�N��U���
�`�
�0��l�C��Y����K+��c�����9�<�9�
�e��(���K����CT�N�����u�f�n�u�w�}�W���Y�����h_�*���
�d�l�i�w�%�(���5����G9��[�����g�
�
� �e�d�(��K�ƨ�D��\�N���u�u�u�u�w�}�WϪ�	����l��hZ�A��u�-�
���$��������_��Y��*���g�l�
�g�b�}��������l�N��U���u�u�u�!�'�l�@�������F���%���:�
�}�d�3�*����H��ƹF�N��U���u�u��6��<��������A��V�����e�g�i�u��>�(�������F��E��AҊ� �g�a�
�d�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߊu�u�x�4�$�:�W�������K��N�����0�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��D���!�0�_�u�w�}�W���Y���N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��1����|�4�1�}�/�)��������V��N�����:�&�
�#��t�^Ϫ����F�N��U���u�4�'�9��2�(���	����lT��h^��*���
�l�u�h�6�/��������\��Z��*���
�
� �f�d��D�ԜY���F�N��Uʴ�'�9�
�:��2���M�ԓ�lW��h��*��u�h�4�'�;���������R��h��*ߊ� �f�b�
�d�W�W���Y���F�N��*������0�:�o�C���I����lT��R�����9�
�:�
�8�-�E���K����lU��B1�G܊�f�_�u�u�w�}�W���Y�Ư�l/��r6��'���8�g�a�0�f�/���L���R��[�����:�%�g�a�e�8�F�������P��UךU���u�u�u�u�w�}����=����a��Z1�C���e�'�2�g�`�a�W���&����\��X��G���g�0�e�d�1��A���	��ƹF�N��U���u�u�9����%�������9��1����a�i�u�'��)�1���5����V��1��D���3�
�c�e�'�f�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠu�u�x�u�$�4�Ϯ�����F�=N��U���6�&�u�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��R��u�=�;�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9�� 1����|�u�=�;�w�}�W���Y���F��d1��<��� �
�d�
�2��@��E�ƫ�C9��h]�*��_�u�u�u�w�}�W���Y����w/��x��D���'�2�f�a�w�`��������9��d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԜY�����^	�����0�&�u�x�w�}�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�F�������F�N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�c�;���P����[��N��U���u�u�u�u�>�����
����A��B��D���g�'�2�a�b�}�JϷ�&����R��d�����0�d�d�g�1��D���	��ƹF�N��U���u�u��6��<��������A�� V��*���
�d�f�i�w���������G��C��*��
�
� �f�g��D�ԜY���F�N��Uʼ�
�!��&��)��������9��E��A��u�h�<�
�#���������F��V��F���
�a�b�%�l�}�W���Y���F���M���2�a�b�u�j�/�ׁ�����9��d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԜY�����^	�����0�&�u�x�w�}�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�F�������F�N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�f�;���P����[��N��U���u�u�u�u�>�0�D�������F���ي� �g�e�
�e�W�W���Y���F�N��#���
�d�'�2�d�e�W��	����9��h��G��
�f�_�u�w�}�W���Y���@��C��E���2�a�e�u�j�.����	�֓�F9��]��G�ߊu�u�u�u�w�}�W�������CS��E��A��u�h�&�9�#�-�E���&����l��=N��U���u�u�u�u�w�8�(���Lǹ��T9��\��Hʦ�9�!�%�a�1��C���	��ƹF�N��U���u�u�8�
�f�/���@�����hV�����a�d�%�n�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװU���x�u�&�<�9�-����
���9F������u�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�_��U���;�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����V��D��\���!�0�_�u�w�}�W���Y���\��Q��*؊�0�
�l�c�k�}��������l ��\�*��_�u�u�u�w�}�W���Y����_T��1����a�u�h�%��1�(�������T��UךU���u�u�u�u�w�}�(���K����A��W�U��%��9�
�g�;�(��J����9F�N��U���u�u�u�8��n�(���&����Z�G1��؊�c�3�
�d�e�-�_������\F��UךU���u�u�u�u�w�}��������9��C1����b�u�h� �3�/����K����l ��\�*��_�u�u�u�w�}�W���Y����A ��@1�����f�b�u�h�"�9�����ԓ�F9�� W��G�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�F܁�
����O�C�����u�u�u�u�w�}�W����ԓ�9��P1�@���h�%��9��k����K�ߓ� ]ǻN��U���u�u�u�u��<�E���Hʹ��T9��X��Hʥ��9�
�
�n�;�(��I����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�}�W��Y����]�������4�
��3�:�}�Ϫ�ӕ��G��V�����x�_�u�u�'��(���&����T��E��Oʥ�:�0�&�}�'�.����Y����`9��ZB�����y�0�<�6�9����Lù��l�N�����u�u�u�u�4�.�W���:����^F��=N��U���u�u�u�=�9�<�(���
�ד�@��S����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t�������R��C��U���%�6�;�!�;�:���P����[��N��U���u�u�u�u�w�}����*����Z�V��!���g�3�8�d�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:��؊�&�
�u�k�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W�������l ��R������&�f�3�:�o�}���Y���F�N�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�����B���F�N��U���u�;�u�3�]�}�W���Y���D����&���!�
�&�
�w�c�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�c�;���s���F�N��U���0�&�_�u�w�}�W���Y���F�V��&���8�i�u�%���܁�
����9F�N��U���u�u�u�;�w�;�}���Y���F�@��U����
�!�
�$��W���s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�B�������F�N��U���u�u�0�&�]�}�W���Y���F�N������3�8�i�w�-�$���ǹ��^9��=N��U���u�u�u�u�w�3�W���s���F�N�����u�%��
�#�����Y���F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����
�&�u�h�6��#���O����lS��N��U���u�u�u�u�2�.�}���Y���F�N��U���4�
��3�:�a�W���*����9��Z1����u�u�u�u�w�}�W���Y����F�N��U���"�0�u�%���ف�
����X�N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���%��
�&�w�`����-����l ��hX�U���u�u�u�u�w�}����s���F�N��U���u�u�4�
��;���Y����g9��1�����_�u�u�u�w�}�W���Y����Z ��N��U���u�u�"�0�w�-�$���Ĺ��^9��
P��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}�W�������F�N��U���u�u�u�u�6��$������R��c1��B���8�c�_�u�w�}�W���Y���V��^�U���u�u�u�u� �8�W���*����9��Z1�H���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W���Y����_��N��U���u�u�u�u�w�}����*����Z�V��!���m�3�8�b�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����g9��1����h�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���e�3�8�l�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:�����3�8�l�h�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�d�1�0�F��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�F߁�
����9F�N��U���u�u�u�;�w�;�}���Y���F�@��U����
�!�d�1�0�F���G���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���;���&�u�h�4��	���&����W��N��U���u�u�u�u�2�.�}���Y���F�N��U���4�
��3�:�a�W���*����W��D��E�ߊu�u�u�u�w�}�W����ƥ�l�N��U���u�"�0�u�'��(���K����lW��
P��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�%���.�W������l��1����n�u�u�u�w�}�W���YӃ��Vl�N��U���u�u�u�u�w�<�(������F��h=����
�&�
�d�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����g9��]�����g�h�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���7����^F���&���!�a�3�8�f�f�W���Y���F�N�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�f�����K���F�N��U���u�0�1�<�l�}�W���Y�����YN��*���&�d�
�&��n�J���Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��h �����i�u�%���)�B�������9F�N��U���u�u�u�9�2�}�W���Y���F�N��U����
�&�u�j�<�(���
����U��]�U���u�u�u�u�w�}������ƹF�N��U���=�;�4�
��.�Fځ�
����[�=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Q����P	��h��F���
�g�h�4��2����¹��O�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���<�u�}�4��2��������F�V�����;�u�0�<�4�3�(���J����CT������!�9�d�e�~�}����Y���F�N��U���u�u�%���.�W������l��1����n�u�u�u�w�}�W���YӃ��Vl�N��U���u�u�u�u�w�<�(������F��h=����
�&�
�a�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����A�	N��U���u�u�u�u�w�}����*����Z�6��-�������u�W�W���Y�Ʃ�WF��D�U���0�1�%�:�2�.�}���Y�ԓ�l ��W�����h�&�1�9�0�>�����ι�@��R
�����;�!�9�d��n�^������]��C��F܊� �a�f�%�~�f�W���?����lU��h�I���!�
�:�<��8��������]��V�����
�#�g�a�d�}�W���������h\�� ��`�%�|�n�w�}�&���&����9��h[�*��i�u�d�u�?�3�_�������9��Q��Lӊ�g�u�u�<�9�9��������_��h_�\ʰ�&�u�e�n�w�}�&���&����U��_��G��u�d�u�=�9�u����۠��U��[��G���u�<�;�1�6�����&����lW��N�����e�n�u�u��3�ށ�����V��h��D��
�g�i�u�#�-�(���H����CT��Y
�����g�3�
�f�g�-�^�ԜY�ƞ�]��h��*���&�g�3�
�f��E��Y۴��T��V�����
�
�d�3��m�(������R��1�����0�
�
� �o�j����s���a��R_�����;�&�g�<��h����N�ӓ�F�F�����d�<�
� �f�m�(������R��1�����0�
�
�d�%�:�D��P���F��Y	��*���
�;�&�g�>����J����[�N��U����;�0�
�;�����K����
W��G\�����}�'�6�;�f�j�ށ�����l��G��U��|�0�&�u�w�}�W���
����^��h��L���%�n�u�u��3�ށ�����V��h��A���
�l�l�%�w�`�_�������Z9��P1�E���;�u�4�2�f�<��������Z9��P1�G���_�u�u�4�0�l��������9��Q��@���%�u�h�_�w�}�W�������l��h�����
�a�m�%�w�5��������WW��h�� ��m�
�g�e�w�}�F�������9F�N��U���
�8�g�
�"�l�Cׁ�J���F��Y	��*���
�;�&�g�:�%�ށ����� 9��R��]���2�d�4�9�8�8�(݁�H����lU��N��ʶ�'�,�d�;�#�4�(���H����CT�=N��U���2�d�4�9�8�8�(݁�����U��_�����h�}�4�2�f�<��������Z9��h_�C���u�;�u�4�%��(���&����lW��1��\�ߊu�u�4�2�f�<��������U��Y��G��u�!�%�
�"�e�F���Y����G��W�� ��b�%�|�_�w�}����H����l	��D1�����b�`�%�u�j��Uϩ�����l4��B��D���
�b�`�%�w�}��������EU��N�����e�n�u�u��3�ށ�����V��h��F��
�g�i�u�f�}����Q����@��hZ�����d�a�h�4��2����������RN��W�ߊu�u�4�2�f�<��������lW��1��U��}�4�2�g�6�1����&¹��U��Y�����;�u�4�2�f�<��������U��\�����_�u�u�4�0�l��������lW��B1�DҊ�g�i�u�d�w�5��������U��]�����u�%�6�;�#�1�Bہ�PӃ��VF�UךU���4�2�d�4�;�'����K����
T��G\��H���4�2�d�4�;�2����&����Q��N��ʴ�
�:�&�
�!��^�ԜY�ƞ�]��h��*���:�
�
�d�1��Nց�J���9F�N��U���g�
�d�3��n�(������	��T��D���<�
� �l�n�-�_���D����F��D��U���u�u�&�9�#�-�F���&����CU��N��'���0�
�9�
�2�2�(݁�&����Q��G]��H�ߊu�u�u�u��o�(�������9�������'�6�;�d�`�4����M�ԓ�N��S��D���0�&�u�u�w�}�Wϭ�����W��B1�Cފ�f�_�u�u�6�:�F�������\��h��L���%�u�h�w�u�*��������lP��B1�@���u�u�%�6�9�)���&����_��^�����u�4�2�d�6�1����
�ғ�F9��_��G��u�d�u�=�9�u�(�������l ��Y�*��h�4�
�:�$��܁�PӃ��VF�UךU���4�2�d�4�;�'����L���� V��h�I���d�u�=�;�������ғ�V��]�Hʴ�
�:�&�
�!��^ϻ�
���]ǻN�����d�4�9�/�%�.����L�֓�F�F�����
�9�
�;�$�l����M�֓�F��EN��*���&�
�#�
�~�W�W�������l0��h��D���
�g�i�u�#�����&����\��_��*���=�}�;�<�9�9����/����V��h�Y���<�!�2�'�"�.����Q���F��G1�*���d�`�
�d�d�p�W������O�UךU���4�2�g��d�;�(��&���F��S1�����#�6�:�}�?�;�(����ι�@��R
�����
�
� �a�b�-�^ê�&����T��B �����}�e�u�u�:��B���&����CW�C����!�u�|�|�~�W�W�������l��h�����3�
�l�
�e�a�W��Y����N��Y	��*���
� �m�f�'�}�W���&¹��l^��h�U���0�w�w�_�w�}����K����l	��D1��ۊ� �l�d�%�w�`�}���Y���a��R\�����;�&�d�3��d�(������	��T��D���<�
� �m�d�-�_���D����F��D��U���u�u�'�#��(�O���	��ƹF��V ��G���9�:�0�
�����Nǹ��Z�=N��U���u�4�2�g�6�1����&����P��G\�����}�'�6�;�f�h����&����l��G��U��|�0�&�u�w�}�W�������U��]����u�u��;�2���������l��h�����b�g�%�u�j�u����K����l	��D1��ۊ�0�
�m�c�/�/��������_��G�U����;�0�
�;�����H����l��B1�LҊ�g�i�u��9�8�(���&����lW��h��D��
�f�-�'�6�����&����O��N��'���0�
�9�
�9�.�D���&����l��S��D���=�;�}�
�2�(����HĹ��lT��1��U���%�6�;�!�;�o�D������D��N��'���0�
�9�
�9�.�C���&����l��S��D���=�;�}�
�2�(��������T��
N��*���&�
�#�
�~�8����I��ƹF��V ��G���9�:�0�
�"�l�Aׁ�K���W�@��U�;�0�
�
��(�F��&�����h��D��
�g�u�9�2��U�ԶY���F��h
��ʴ�&�2�u�'�4�.�Y��s���R��X �����2�
�'�6�m�-����
ۇ��@��CB�����2�6�0�
��.�F������R��RB�����2�6�0�
��.�Fځ�
����F��^����� �f�`�
�e�W�W�������F�N�����}�;�!�}�'�>��������lW������!�|�4�1��-��������Z��S�����2�6�0�
��.�F������	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��@���8�d�|�4�3�3��������]��B1�@ڊ�g�h�4�
�8�.�(���&���O��_�����u�u�u�u�w�-����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�:�0�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�4�
�3�8�����Ƽ�\��D@��X���u�4�
�1�2�<����&����\��E�����%�&�4�!�w�-��������`2��C_�����|�u�u�7�0�3�W���Y����UF�Y��]���6�;�!�9�0�>�F������R��N�����%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�t�W������F�N��Uʴ�
�1�0�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��[��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������,�4�&�2�w�/����W���F�V�����
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	���&����R�R�����
� �f�`��o�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�`�1�0�F�������\�R�����
� �f�`��o�JϿ�&����G9��1�\���!�0�u�u�w�}�W���YӇ��A��NN�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����F��N�����u�'�6�&�y�p�}���Y����V��Y1�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�h����H����K��X �����a�e�%�y�6�/��������\��Z��*���
�
�0�
�n�q��������lV��E�����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���4�1�;�!��%�������� R��h�Hʴ�
�:�&�
�!��^���Y����l�N��U���u�4�
�0�"�3�G��Y����_��X�����g�a�g�0�g�k����K����F�N�����u�u�u�u�w�}�WϿ�&����A��R�����0� �;�e�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����
�u�&�<�9�-����
���9F������'�
�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
����U��Z����6�;�
� �d�h�(��Y����_��X�����g�a�g�0�f�k����K���R��R�����%�0�|�u�w�?����Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�a�w�3�W���Qۃ��G��S1��*��e�%�u�u�'�>�����ד�O����ߊu�u�u�u�w�}��������F���*����'��:��m�(݁�&¹��A��X����u�u�u�9�2�W�W���Y���F��h�� ���d�i�u�%�%�)����&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�0� �9�o�����Ƽ�\��D@��X���u�4�
�0�"�3�E���
����C��T�����&�}�%�6�{�<�(���&����l5��D�*���
�a�u�-�#�2����&����l����<�����!�'��n�(���&����^�������'�
�
�'�0�W�W�������F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�`�3�:�l�^Ͽ�ӈ��N��^����� �f�`�
�e�`��������_��G��\ʡ�0�u�u�u�w�}�W�������G��h\��Hʶ�
�����8���M����l��h\�N���u�u�u�0�$�}�W���Y���F��G1�����
�u�h�4��8����K����T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�'�!�%��W�������A	��D�X�ߊu�u�%�'�#�/�(܁�
����l��TN����0�&�4�
�2�}��������B9��h��@���8�d�y�0�>�>��������9��N��*������0�:�o�C���H����lT��N��*��� �;�f�%�2�t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��C����Ƣ�GN��O�����3�
�a�e�'�}�W�������l
��h^��\���=�;�_�u�w�}�W���Y����V��Y1�I���9�����)����Jǹ��9��P1�@�ߊu�u�u�u�;�8�}���Y���F�V�����;�f�i�u�'�/����&����V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�4�
�0�"�3�CϿ�
����C��R��U���u�u�4�
�2�(��������]9��X��U���6�&�}�%�4�q��������V��c1��Dߊ�&�
�a�u�/�)��������V��B��������!�%��Dف�&ù��T9�� B�����!�'�
�
�%�:�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�`�1�0�F�������\�R�����
� �f�`��o�JϿ�&����G9��1�\���!�0�u�u�w�}�W���YӇ��A��E ��U��6�
��������K�Г�lV��R	��B��u�u�u�u�2�.�W���Y���F������'�
�u�h�6������ғ�A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�%�'�#�/�(���
������T��[���_�u�u�%�%�)����&����T��E��Oʥ�:�0�&�4��8�W���
����@��d:�����3�8�d�y�2�4����&����S��G\��������2�0�E����ד�V��Z����0� �;�`�'�8�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(��Y����]	�������1�3�
�a�g�-�W���	����@��A_��\���u�=�;�_�w�}�W���Y�ƭ�l��B��@��u�9��������&����V9��E��G��_�u�u�u�w�1��ԜY���F�N��*��� �;�`�i�w�-��������C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�4�
�>�����J�ƭ�@�������{�x�_�u�w�-�������� U��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��F���h�}�%�6�9�)����H����C9��h��]���:�;�:�m�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����L�ƭ�@�������{�x�_�u�w�-��������Q��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��@���h�}�%�6�9�)����H����C9��h��]���:�;�:�l�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����N�ƭ�@�������{�x�_�u�w�-��������Q��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��B���h�}�%�6�9�)����H����C9��h��]��1�"�!�u�g�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����d�1�"�!�w�l�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������
T��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��^�*���<�;�%�:�w�}����
�έ�l%��Q�����u�0�<�_�w�}�W���Y���F��h��*���
�e�g�i�w�<�(���
����9��
N��*���3�8�d�1� �)�W���B����������n�_�u�u�z�}��������lT��N�����u�'�6�&�y�p�}���Y����Z��S
��D���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�g�e�w�`�_�������l
��h_��U����
�&�}�w�2����K����F�R �����0�&�_�_�w�}�ZϿ�&����Q��_�U���<�;�%�:�2�.�W��Y����C9��P1����e�
�&�<�9�-����Y����V��V��&���8�_�u�u�2�4�}���Y���F�N�����<�
�1�
�f�e�K�������]��[��D��4�
��3�:�n��������]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��D���4�&�2�u�%�>���T���F��h��*���
�d�`�4�$�:�(�������A	��D�����
�&�|�u�w�?����Y���F�N��U���%�&�2�7�3�o�F���D�έ�l��D��ۊ�u�u�%���.�_�������R�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����g�u�&�<�9�-����
���9F������7�1�g�g��.����	����	F��X��´�
��3�8�]�}�W������F�N��U���u�4�
�<��9�(��J�����T�����d�d�h�4������Lӂ��]��G����u�;�u�'�4�.�L�ԶY���F��h��*���
�a�u�&�>�3�������KǻN�����2�7�1�g�n�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���@�����T�����d�d�h�4������H�ƨ�D��_�\�ߊu�u�;�u�%�>���s���K�V�����1�
�c�u�$�4�Ϯ�����F�=N��U���&�2�7�1�e�l��������\������}�%��
�$�t�W�������9F�N��U���u�u�u�%�$�:����K���F��G1�����9�d�d�h�6��$�������W	��C��F���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�b�`�<����Y����V��C�U���4�
�<�
�3��@�������]9��X��U���6�&�}�%�$�:����&����GW��Q��D���0�<�6�;��(�D��&���F�U�����u�u�u�u�w�}�WϿ�&����Q��Y�U��}�4�
�:�$�����&���R��^	������
�!�`�1�0�F������V��T��*���f�`�
�g�j�<�(���
����9��UךU���;�u�'�6�$�f�}���Y���R��^	�����b�u�&�<�9�-����
���9F������7�1�g�b�6�.���������T��]����
�&�|�w�}�������F�N��U���u�%�&�2�5�9�E��E����C9��Y�����d�h�4�
��;���Y����G	�G����u�;�u�'�4�.�L�ԶY���F��h��*���
�f�4�&�0�}����
���l�N��*���
�1�
�f�6�.���������T��]����
�&�|�w�}�������F�N��U���u�%�&�2�5�9�D���D�έ�l%��Q��Eʱ�"�!�u�|�j�<�(���
����9��d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����u�&�<�;�'�2����Y��ƹF��G1�����1�c�
�&�>�3����Y�Ƽ�\��DF��*���3�8�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��d�K�������]��[��D��4�
��3�:�k��������]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��Dʴ�&�2�u�'�4�.�Y��s���R��^	�����d�4�&�2��/���	����@��G1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�m�w�`�_�������l
��h_��U����
�&�}�w�2����N����F�R �����0�&�_�_�w�}�ZϿ�&����P��h=����
�&�
�u�$�4�Ϯ�����F�=N��U���&�2�6�0��	���&����
9��D��*���6�o�%�:�2�.��������W9�� GךU���0�<�_�u�w�}�W���Q����Z��S
��@���!�0�u�u�w�}�W���YӇ��@��T��*���&�d�
�&��}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�m����@���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���d�
�&�
�g�<����Y����V��C�U���4�
�<�
�$�,�$����ד�@��1�����
�'�6�o�'�2��������T9��S1�B�ߊu�u�0�<�]�}�W���Y���R��^	�����b�|�!�0�w�}�W���Y�����D�����
��&�d��.�(��E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	���&����V�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����D�����
��&�d��.�(������]F��X�����x�u�u�4��4�(�������@��h��*���4�&�2�
�%�>�MϮ�������D�����d�b�_�u�w�8��ԜY���F��F��*���
�1�
�l�~�)����Y���F�N�����2�6�0�
��.�F݁�
����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����9��Z1�U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C�����2�6�0�
��.�F܁�
������^	�����0�&�u�x�w�}��������V��c1��Dي�&�
�g�4�$�:�(�������A	��D�����2�7�1�g�n�W�W�������F�N�����4�
�<�
�3��C�������9F�N��U���u�%�&�2�4�8�(���
����U��\��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��C_�����d�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
����U��]�����;�%�:�0�$�}�Z���YӇ��@��T��*���&�d�
�&��n��������\������}�%�&�2�5�9�E��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���a�3�8�d�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�.��������l��1����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�f�����M����Z��G��U���'�6�&�}�'�.��������l�N�����u�u�u�u�>�}��������W9�� G�����_�u�u�u�w�}�W���
����@��d:�����3�8�d�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�`�1�0�F���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����@��d:��ۊ�&�
�u�&�>�3�������KǻN�����2�6�0�
��.�F����֓�@��Y1�����u�'�6�&��-�������� OǻN�����_�u�u�u�w�;�_���
����W��G�����_�u�u�u�w�}�W���
����@��d:��ۊ�&�
�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��C\�����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�e�;��������]9��X��U���6�&�}�%�$�:����K����9F����ߊu�u�u�u�1�u��������lT��G�����_�u�u�u�w�}�W���
����@��d:��؊�&�
�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��C]�����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�d�;��������]9��X��U���6�&�}�%�$�:����K����9F����ߊu�u�u�u�1�u��������lT��G�����_�u�u�u�w�}�W���
����@��d:��ي�&�
�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��CZ�����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�c�;��������]9��X��U���6�&�}�%�$�:����K����9F����ߊu�u�u�u�1�u��������lT��G�����_�u�u�u�w�}�W���
����@��d:��ފ�&�
�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��C[�����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�b�;��������]9��X��U���6�&�}�%�$�:����K����9F����ߊu�u�u�u�1�u��������lT��G�����_�u�u�u�w�}�W���
����@��d:��ߊ�&�
�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��CX�����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�a�;��������]9��X��U���6�&�}�%�$�:����K����9F����ߊu�u�u�u�1�u��������lT��G�����_�u�u�u�w�}�W���
����@��d:��܊�&�
�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��CY�����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�`�;��������]9��X��U���6�&�}�%�$�:����O��ƹF��R	�����u�u�u�3��-��������
O��_�����u�u�u�u�w�-��������`2��CY�����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����G^��D��U���<�;�%�:�2�.�W��Y����C9��P1������&�m�3�:�j��������\������}�%�&�2�5�9�O���Y����V��=N��U���u�3�}�%�$�:����A����[��=N��U���u�u�u�%�$�:����&����G^��D��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}��������B9��h��*���
�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
�ߓ�@�������%�:�0�&�w�p�W�������T9��R��!���l�3�8�m�6�.���������T��]���&�2�7�1�f�n�}���Y����]l�N��Uʼ�u�4�
�<��9�(��PӒ��]FǻN��U���u�u�%�&�0�>����-����l ��hV��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��CW�����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǻN��U���'�
�!��%�����Iǹ��V9��Q��@���%�u�h�&�3�1��������AN��D��]���;�1�!�%�f�i����L�֓�O�G����u�4�'�9��2�(���	����lV��h_�� ��m�
�g�i�w�)�(�������P�������4�'�9�
�8�����K�ғ�l��h��F��
�d�u�u�>�3�Ƿ�&����9��h<�����;�
�:�'�2�o����L�ѓ� O�=N��U���
�!��'��2�(��&����9��Q��C���%�u�h�_�w�}�W�������v>��e����c�0�e�'�0�o�@ϩ�����V
��Z�*���f�e�
�g�g�}�W��PӃ��VFǻN��U���'�
�!��%�����Iǹ��V9��Q��@���%�n�u�u�6�/��������\��Z��*���
�
� �f�f��D��Y���F���*����'��:��m�(߁�&ù��lU��1��U���;�}�0�
�:�e����L�֓�N��S��D���0�&�u�u�w�}�WϽ�&����k'��C��*��
�
�
�0��e�L���YӇ��l
��q��9���
�e�
�
���(���J����CU�
NךU���u�u�9����%�������9��1����m�"�0�u�$�1����I���� P��h�E���u�d�|�0�$�}�W���Y����A��C1�����:�
�e�
���(݁�����9��d��Uʴ�'�9�
�:��2���M�ԓ�lV��h��F��
�f�i�u�w�}�W�������G9��E1�����e�
�
�
��(�D��&����[����*���d�
� �f�g��E��Y���O��[�����u�u�u�'��)�1���5����V��1��E���'�2�g�l�]�}�W���&����\��X��G���g�0�e�3��h�A���Y���F�N���������2�0�E����֓�V�� Y�����}�0�
�8�o�;�(��I����O�I�\ʰ�&�u�u�u�w�}��������A9��X��Eފ�
�
�
� �d�e�(��s���R��[�����:�%�g�a�e�8�F�������V��N�U���u�u�u�6���2���+����lT��h��*���
�a�u�=�9�u��������U��^�����|�h�r�r�w�1��ԜY���F��E1��*���
�:�%�g�c�o��������T��UךU���'�
�!��%�����Iǹ��V9��1��*��m�%�u�h�]�}�W���Y����_��X�����g�a�e�0�f�;�(��M����D��F�����%�
� �f�n��E��Y���O��[�����u�u�u�9���/�������U��R1�����g�`�_�u�w�/�(���?����\	��^��G���d�f�3�
�a�k����D���F�N��*������0�:�o�C���H����lT�������0�
�8�d��(�D��&���F�_��U���0�_�u�u�w�}��������l*��G1�A���0�d�g�3��k�O���B�����h��3����:�
�e���(ށ�&����Q��G]��H�ߊu�u�u�u�%���������C9��1�����3�
�`�a�'�}����Q����G��1��*��a�%�}�|�j�z�P������F�N�����9�
�:�
�8�-�E���K����lP��R	��C��u�u�4�'�;���������R��h��*���f�a�
�f�k�}�W���Y����_9��s+��'���'�
�f�
������M�ƻ�V�D�����
� �f�l��o�G���Y�����RNךU���u�u�'�
�#���������9��R1�����`�a�%�n�w�}����&����|��p������
�$�4�����L¹��Z���*��
� �g�a��n��������]��[��D��u�u�7�:���G���&����G��x�����
�
� �g�n��E��Yے��lW��h��*��`�-�'�4��2����¹��l�N������,� �
�%�<��������R
��h��G��
�g�i�u�"�)����J�ѓ�F��EN��*���&�
�#�
�~�W�W�������VW��h
�����;�<�
� �f�n�(��E����V��P �����3�
�b�d�'�}��������W9��R��*���3�
�b�d�'�t�}���Y����A��_�����2�;�<�3��m�O���Y���]��^	�����0�
�l�d�6�9��������]��1�����l�a�%�|�]�}�W�������W��1��*��a�%�u�h��/����H�ד�V��P��ۊ� �d�f�
�e�%�Ͽ�&����G9��1�N���u�7�8�'�2�o�(������� 9��R��]���0�2�d�d�3�0����&����lT��1��U���u�%�6�;�#�1�F��B�����R��D���<�
� �d�c��E��Yۅ��A��h ��*���3�
�b�c�'�}�ό�����R
��X ��*ۊ�:�
�d�3��j�E���P���F��Z����
�
� �d�g��E��Yۅ��A��h ��*��� �d�l�
�e�2�W����ԓ�_
��Y��D���!�<�3�
�b�e����s���Q��E	��*���d�b�
�g�k�}����H����^��h����'�0�2�d�f�9��������l ��V�*��n�u�u�7�:�/��������T��^_�� ��b�
�g�i�w�3� ������� 9��h\�F���u�;�u�0�2�8�(���
�ԓ�F9��V��F��u�u�7�8�%�8�G�������]9��h��F���
�g�i�u�9�*��������U��X�����;�u�0�0�2�����J���� W��h�N���u�7�8�'�2�m��������Z9��h\�B���u�h�}�<�9�4�(���K����CU��Y
�����2�7�!�g�1��F���	����F�U�����3�
�e�f�'�}�J����ӓ�F9��Y��Gʺ�u�'�0�2�f�l��������Z9��h\�M���|�_�u�u�%�8����H����^��h�I���;�"�<�;�>��(���H����CU��EN�����1�/�'�&�g�3����&����W��G\����u�'�0�2��o����K�ӓ�F�F�����;�<�
�
�"�o�Nց�JӉ��C9��C1�����g�l�%�|�]�}�W�������ZU��B1�@܊�g�i�u�;� �4����&����lT��1��U���%�;�!�<��(�E��&���9F������
�a�3�
�f�h����D�΢�D��Y��*ފ� �f�c�
�d�2�W�������l ��_�*��n�u�u�7�:�/��������T��N�U»�"�<�;�<��8�(��HӉ��W��C�����&�e�;�!�>�;�(��N����l�N�����0�<�<�
�"�l�Bف�K�����R�����
� �d�`��o��������\��h��D��
�g�n�u�w�?��������9��h\�L���u�h�}�;�2�;����&���� _�������3�:�
�
�2��N��B�����R��*���f�3�
�l�a�-�W��Q����A ��@1�����l�d�%�u�%�2��������U��X�����_�u�u�'�2�:�(���M���� W��h�I��� �1�'�9� �i����H�֓�F�������"�a�3�
�f�k����s���Q��E	�����3�
�e�`�'�}�J�������_	��Q��E���%�u�'�:�2�;��������9��UךU���4�'�
�
�"�o�F؁�K�����h_�*���
�e�d�4�3�)���&����
W��G\����u�4�'�
��l����N�ӓ�F�F�����%�g�3�
�a�d�����Ƹ�CQ��B1�Lӊ�g�n�u�u�4�/��������U��h�I���&�9�!�%�f�;�(��J����R��C��*���d�a�
�g�l�}�WϽ�����l��h�����b�c�%�u�j�u�������� W��N��U���
�g�
� �f�h�(��B�����E��*���
�
� �d�n��E��Yے�� 9��h_�C���u�'�!�%�a����LŹ��]ǻN�����
�
� �f�`��E��Yے��lW��h��*��a�4�1�!�'�d�(���J����CT�=N��U���'�
� �g�f��E��Yے��lW��h��G��
�f�4�1�#�-�@ځ�����9��UךU���0�0�0�
�9�.�G���&����^��G\��H���0�0�0�
�9�.�F���&����l��X�����8�a�
� �f�j�(��B�����R��*���&�e�<�3��d�C���Y���W��C�����
�0�
�l�a�2�W���&����9��h_�L���|�_�u�u�2�8��������l ��Y�*��i�u�u�u�w�}�%���¹��_9��R��*���
�d�3�
�`�n�������Q��E	��Gي�d�3�
�b�`�-�_���D����F��D��U���u�u�%�d�g�4�(���&����l�N�����1�:�0�
��(�E��&���FǻN��U���
�d�<�
�"�o�D܁�Kӑ��]F��V��*ۊ� �g�d�
�e�m�W���H����_��=N��U���u�4�2�d�6�1����&ƹ��T9��_�U���1�9�!�1�8�8�(܁�����9��R�����u�u�u�
�f�4�(���J����CT��_��]���'�
�
� �d�j�(��I���W����ߊu�u�u�u�6�:�F�������@9��Q��E���%�n�u�u�3�1��������U��]�����h�_�u�u�w�}����H����l	��D1�����<�3�
�c�g�-�W����ή�^��R_�*��� �d�e�
�e�m�W���H����_��=N��U���u�
�g�
��(�F��&����F�S�����/�'�&�e�9�)�ށ�����9��R��]���
�l�'�2�d�k�W���Y����G��M�����;�!�3�
�o�m����s���W��C�����&�e�;�!�>�;�(��N����[�C��G؊�0�
�l�m�6�9��������V��h ��*���d�l�
�g�l�}�WϺ�����l��X��*���d�d�
�f�k�}�W���Y����R��1�����0�
�
�d�%�:�D��Y����N��E��D���
� �d�e��o�G���Y�����RNךU���u�u�4�2�f�<��������l��E��F��n�u�u�1�;�)��������l��h��D��
�g�i�u�3�1��������lW��B1�Dӊ�f�-�'�4��2����¹��l�N�����1�/�'�&�e�;�(��H����[�D�����3�
�d�d�'�}��������A��Q��G���%�|�_�u�w�8����&����@9��Q��L���%�u�h�_�w�}�W�������l��h�����'�2�a�m�w�5��������9��h\�B���}�|�h�r�p�}����s���F�e��ۊ�9�
�0�:������I����F�S�����/�'�&�a�1��G���	���l�N��Uʇ�;�0�
�9��3��������P��N�����6�'�,�g�1��G���	����[�I�����u�u�u�u�w�����&����I��D1�����e�d�%�n�w�}��������V��h��D��
�f�i�u�w�}�W���+����9��[1�����
�
�0�
�n�h� ���Yۅ��A��h�����l�`�e�u�w�l�^ϻ�
��ƹF�N�����d�4�9�/�%�.�E�������
U��=N��U���0�0�
�0�8���������9��R��]���0�0�
�0�8����Mǹ���������!�9�d�d�l�}�Wϻ�����W9��h]�E���u�h�w�w� �8�WǷ�&����\��X�����2�f�e�h�6�����&���� O��[��W���_�u�u�-���(���M�ѓ�F���*���<�
�0�!�%�.����Q����\��h��G���d�u�u�<�9�9����JŹ��lR��h�\�ߊu�u�-�
��(�D���	�����h�����0�!�'�&�0�8�_�������l
��1��D���u�<�;�1�#�-�E���&����CW�d��Uʰ�%�!�%��f�;�(��&���F��R	��*ۊ� �a�b�%��o��������]ǻN�����8�
�
� �d�h����Dӏ��T9��Q��Fӊ�d�c�u�:�9�2�B���s���U��v,��:����&�9�!��<����N�ד�F9��\��F��u�u�u�u�w�-�!���&�Г�V��Z����u�!�%�b��(�E��&���F�_��U���0�_�u�u�w�}����;����G9��D�����4� �
�b�$�;�(��N����9F���*���-� �
�7�8�(��������9��Q��F���%�u�h�&�3�1��������AN��D�����%�6�;�!�;�o�(���Tӓ��Z��SF��#���
�c�'�2�d�i�^��Y����K��u=�� ���7�:� �0��1���&¹��lT��1��U��_�u�u�u�w�����M¹��lT��1��U���;�}�8�
�`�;�(��N����O�I�\ʰ�&�u�u�u�w�}����8����F��U�� ����9�0�l�����O����l�N�������!��$�1��������
_��h��G��
�g�i�u�#�����&����\��Y�����4�
�:�&��+�C��Y�ƹ�@��R
��*���g�a�
� �e�n�(��P���F��G1�����0�8�a�b��;�(��M����[��C
�����
�0�!�'�"�.����Q����\��h��@��u�u�;�<�9�9��������G��h[�*��� �g�l�
�f�t�}���Y����]	��h�����d��3�
�b�n����Dӕ��l
��^�����'� �&�2�2�u��������ET��G��U���<�;�1�3�'�3��������P��h��G��
�d�|�_�w�}�W�������W��R��@����3�
�`�g�-�W��
����\��h�����'�&�/�}�>�3�Ǯ�/����W��R	��L��y�`�|�_�w�}�W�������\��C��*��
�
� �g�n��F��Y����_	��T1�����}�0�<�0�$�:����&����lW��E��F��|�g�|�n�]�}�W���&����9��1�����l�c�%�u�j�W�W���Y�Ƽ�e��h_�����3�
�m�e�'�}����Q����G��1��*��d�%�}�|�j�z�P������F�N�����!�%�c�3��d�E���B��� ��h��9��� �
� �!�'�$�F���/����P��h�I���8�
�m�3��k�B���Q���W��X����n�u�u�3�'�%�"���6����F
��G��D����3�
�c�n�-�W������l ��X�*��_�u�u�-���;�������_��[��Gފ�
� �g�m��o�K�������T��A�����0�<�0� �$�:��������T��A�����<�;�1�3�'�%�"���6����F
��G��D����3�
�c�n�-�^���
����WN��G1�� ����!��9�>�1�(��&����lT��1��\���u�b�|�_�w�}����4����|��z�����
�g�
�
�"�o�Nց�I���G��V�� ��m�
�d�f�w�}�W������]ǻN�������,� ��(���� ����l0��B1�Lӊ�d�i�u�
�����Nƹ��l�N����� ���!��1����&����e9��h\�L���u�h�&�1�;�:��������A��M�����;�1�&�1�;�:��������@��R
�������,� ��(���� ����l0��B1�Lӊ�e�u�u�<�9�9��������J)��h#�����,�d�b��1��A���	���F��G����u�x�2�%�1��Eށ�Ӈ��Z��G�����u�x�u�u�0�-����K¹��l��^	�����u�u�'�6�$�u�������R��^	������
�!�
�$��[Ͽ�&���R��^	������
�!�
�$��[Ͽ�&����P��h=�����3�8�d�u�'�.��������l��h��*���4�
�<�
�$�,�$���ǹ��^9�������6�0�
��$�h����M�ƭ�l��h�����
�!�
�&��t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�}�%�6�9�)���������D�����
��&�d�1�0�G����Ƣ�GN��G1�����h�4�
�:�$�����&���	�������!�9�2�6�f�`��������V��c1��B���8�c�u�'��-��������Z��S�����2�6�0�
��.�E������\�V�����
�:�<�
�w�}��������B9��h��*���
�|�:�u�6�����&����P9��
N��*���
�&�$���)�(���&����AF��G1�����9�2�6�d�j�<�(���&����l5��D�����a�u�'�}�'�>��������lW������6�0�
��$�k����L�����YNךU���u�u�u�u�%����H����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�2�%�3��o�(���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϹ�	���� T��T�����;�%�:�0�$�}�Z���YӁ��l ��\�����&�<�;�%�8�}�W�������R��C��Yʴ�
�<�
�&�&��(���&����J��G1��Yʴ�
�<�
�&�&��(���&����J��G1�����0�
��&�e�;���Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�����f�u�%�&�0�>����-����l ��hZ����<�
�&�$���ف�
����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V �����}�%�&�4�#�`��������_	��T1�\���'�}�%�6�9�)���������D�����
��&�b�1�0�A����έ�l��D�����
�u�u�%�$�:����&����GT��D��\ʺ�u�4�
�:�$�����&���R��^	������
�!�
�$��^ϱ�Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���}�%�6�;�#�1����H����C9��P1������&�`�3�:�i�W���Q����\��h�����u�u�%�&�0�>����-����l ��h[��\���=�;�_�u�w�}�W���Y����U��Y����u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}��������9��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��ԶY����9��h-�����'�6� �0�f�l�E���&����l��S��U���u�u�;�"�2�l�(���J����CU��_��]���6�;�`�3��n�F���Q���A��N�����u�u�u�u�9�*���&���� R��G]�U���<�
�!��$���������Q��Q��G���%�u�h�&�3�1��������AN��P ��]���6�
�4�0��/��������l ��\�*��u�u�<�;�3�-�!���&����l��hZ�C���_�u�u��4�����*����G��h_�*ۊ� �f�e�
�d�a�W���Y�����d��@���
�f�m�%�w�5��������WS��B1�Cۊ�g�e�u�u�f�t����Y���F� ��&���a�3�
�f�f�-�L���Y�����T������'�6� �2�l�O���&����l��S�����:�<�
�0�#�/�����ο�T����*���3�
�g�c�'�t�D���B���F��h��6���
�!� �!�%��Oځ�&����U��G]��H�ߊu�u�u�u�2���������_��N�����:�
�:�1��(�D��&���F�_��U���0�_�u�u�w�}�����ѓ�F9��\��F�ߊu�u��6��<��������A��[�� ��a�
�g�i�w�)�(�������P�������1�<�
�!��.�(�������V9��1��*��e�%�|�x�"�.����Q����_T��1����`�|�n�u�w�4�(���?����\	��W�����a�c�%�u�j�.��������V��EF�����0�}��9��2�(���	����V��^��^ʠ�&�2�0�}�'�>�����ԓ�O��N�����:�0�!�'��n�(���J����CT�
N�����2�6�#�6�8�u��������^��h��F��
�g�u�u�9�4����	����9��W�����d�c�|�_�w�}�;����ד�]9��Y	������0�6�
��(�D��&���FǻN��U���%�6�;�!�;�n�(������@��C��*���f�`�
�g�g�}�W��PӃ��VFǻN��U���0�
�8�a�1��B���	��ƹF��{1�� ��� �
�e�
�"�n�Aځ�K���@��[�����6�:�}�;�>�3�Ƿ�&����\��N� ���2�0�}��#�/�F���&����V9��S1�����
�
� �f�b��D���s���Z��1��*��
�g�i�u�f�}����Q����V��Z��G݊� �b�`�%�~�a�����έ�l��D��Ҋ�|�u�9�0�u��}���Y����9��hY�*��i�u�d�u�?�3�_�������^��V�� ��d�%�|�k�$�:����	����@��A_��E���0�&�u�e�l�}�WϷ�����]	��Q��A���%�u�h�}�4�-�(���K����CT��X�����;�!�9�d�f�f�W�������l ��Z�*��i�u�d�u�?�3�_���&����U��W�����u�%�6�;�#�1�E��Y����D��d��Uʼ�8�
� �a�f�-�W��[����[�������!�%�b�
�"�i�F���P����Z��SF��*���&�
�#�d�g�t����Y���9F���%���:�
�
��;���������l ��[�*��i�u�u�u�w�}��������lR��_��]���
�e�
� �d�j�(��I���W����ߊu�u�u�u��1�(���&����lT��h��F��
�`�_�u�w�/����H����T��G_��Hʱ�4�&�2�
��(�D���	��ƹF��E��#���
�f�
�d�k�}�(�������F9��1��N���u�<�;�2�f�;�(��&���F��R	��*ۊ� �a�b�%��n��������]ǻN��1���3�
�f�
�f�a�W���&�ԓ�F9��1��]���u�u�:�;�8�m�L���Yӊ��U��_�����h�!�%�g��(�F��&���K�
�����e�n�u�u�:�3�!������� T��N�U���
�:�<�
�2�)�ǫ�
����WN��h�����#�a�e�u�w�3����ۖ��V��C1�����e�m�%�|�l�}�Wϳ�����l ��Y�����h�&�1�9�0�>�����ι�@��R
�����;�!�9�`��t�Zϫ�
����WN��e�����
� �a�`�'�t�L���YӋ��l0��h��A���%�u�h�_�w�}�W������� 9��hZ�*��"�0�u�<�9�:�F���&����CU�N��R��u�9�0�_�w�}�W���&����_��h��A���%�n�u�u�:�3�!���&����l��S��U���u�u�8�;��l����I�ԓ�F��R �����2�'�2�f�b�u�^��^���V
��d��U���u�%��&�;��(���H����CW��N�����0�d�
� �d�i�(��E��ƹF�N��9���
�4�0��%�>����H�ד�F9��^��Gʢ�0�u�&�9�#�-�C�������N��S��D���0�&�u�u�w�}�WϷ�&����R��d�����0�d�`�3��o�B���B�����d��D���
�f�f�%�w�`�}���Y���]��R�����f�m�%�u�?�3�_�������l ��]�*��e�u�u�d�~�8����Y���F��R��Ҋ� �f�f�
�d�W�W�������T��B1�Bߊ�f�i�u�u�w�}�WϷ�&����R��d�����0�d�`�3��o�B���Y����N��[1�����3�
�f�g�'�u�^��^���V
��d��U���u�<�
�!��.�(�������V9��1��*��e�%�n�u�w�3� ���H����lU��1��U��_�u�u�u�w���������G��C��*��
� �f�f��l� ���Yە��l��W�� ��b�
�g�e�w�}�F�������9F�N��U���6�
�4�0��/��������l ��\�*��_�u�u�0��1�C���&����l��S��U���u�u�<�
�#���������F��Y�����g�c�%�u�?�3�_���&����9��P1�D���|�h�r�r�w�1��ԜY���F��h��6���
�!� �!�%��@ށ�����9��d��Uʻ�"�0�d�
�"�n�Nׁ�J���9F�N��U����9�g�3��n�B���Y����N��h��ي� �f�g�
�e�m�W���H����_��=N��U���u�0��9�d�;�(��J����9F� ��&���c�3�
�a�c�-�W��s���F�^"�����&�
�!� �#�/�(��&����U��G_�����}�0�
�8�a����H����V�
N��R���9�0�_�u�w�}�W�������@��C�����
�m�
� �d�i�(��s���]��R�*���f�g�
�f�k�}�W���Y����9��h-�����'�6� �0�f�h����K�ӓ�F��R �����!�%�a�'�0�i�F���P���A�R��U���u�u�u�<��)�4���&����P��R1�M���
�g�c�%�l�}�Wϰ�����9��h]�L���u�h�_�u�w�}�W���*����l ��Z�*��"�0�u�:��2�܁�����9��^��H��r�u�9�0�]�}�W���Y����G9��D�����!�'�
�b��(�D��&����F�Y�����3�
�`�d�'�}�J�ԜY���F��G1�����0�8�`�d��;�(��J����D��F��*���1�3�
�`�a�-�_���D����F��D��U���u�u�;�"�2����Kù��l�N�����g�3�
�c�g�-�W��s���F�Q�����
�0�8�`�g�����M�ד�F��R �����m�
�0�
�n�n�G���Y�����RNךU���u�u�-�
�8�8����&����e9��h\�F���n�u�u�u�w�3� ���J�ޓ�R��Q��@���%�u�h�&�3�1��������AN��D��]���;�1�;�"�2�d����L�ד� O�G����u�;�"�0�d�;�(��J����[�N��U���3�%�;�1��8���N����F9��Z��Gʢ�0�u�&�9�#�-�C�������N��S��D���0�&�u�u�w�}�Wϸ�	����V9��E��Eۊ�
� �g�e��o�}���Y����V
��Q��@���%�u�h�_�w�}�W�������W��R��@����3�
�`�g�-�W����θ�C9��h��*��f�e�u�u�f�t����Y���F���*���0�!�'�
�n��(���K����CT��N�����0�`�3�
�b�j����D���F�N�����f�3�
�`�d�-�W����Σ�l��S1��*���c�%�}�|�j�z�P������F�N�����;�1�
�0�:�h�G�������
W��UךU���0��9�
�"�o�G؁�J���9F�N��U����9�a�
�6�)����L�Г�F��R �����:�1�3�
�b�k����P���A�R��U���u�u�u�3�'�3��������
Q��h��G��
�g�_�u�w�8�$���&���� W��G]��H�ߊu�u�u�u��>�(�������F��E��Bۊ� �f�a�
�e�*����
����^��h��F��
�g�e�u�w�l�^ϻ�
��ƹF�N��9���
�4�0��%�>����H�ޓ�F9��X��D�ߊu�u�0��;����J����Z�=N��U���u��6�
�6�8�$�������lW��h��F��
�g�"�0�w�.����	�ߓ�F9�� X��G��u�u�d�|�2�.�W���Y�����T������'�6� �2�l�O���&����l��=N��U����9�
� �e�d�(��E��ƹF�N��*���g�a�
�0��d�Eϩ�����V
��Z�*���
�e�g�e�w�}�F�������9F�N��U���4�g�d�
�2��N��s���]��R�� ��g�
�f�i�w�}�W���YӀ��l��R1�����e�
�
� �e�m�(��������h��@ڊ�0�
�e�e�g�}�W��PӃ��VFǻN��U���-�
�:�0�#�/�(��&����lT��1��N���u�;�"�<�9�4�(ށ�����9��R�����9�
�l�3��k�O���Q����\��XN�\�ߊu�u�0�&�0�?��������
_��N�U���4�g�f�
�"�o�N܁�K����W	��C��F��u�u�;�"�>�3����&����
V��G]��Hʥ��9�
�d�1��O���	������Y��F���_�u�u�0�$�:����M���� V��h�I���
�4�g�`��(�D��&���F��@ ��U��n�u�u�;�#�>��������S��N�U»�"�<�;�<�����@ʹ��	��G1�����
�a�;�!�1��E���	����F�X�����d�
�d�3��j�(��E����^��1��*��
�g�4�1�%�+�(���A�ד�O��N�����:�1�d�
��(�F��&���F��Z��B���
�a�e�%�w�3�W���H����R��h�N���u�:�
�:�3�l�(�������
9��R��]���
�a�3�
�a��EϿ�Ӕ��9��hV�*��n�u�u�:��2���&����lW��1��U��}�8�
�b�1��C���	�ƭ�WF��A1��*��a�%�|�_�w�}�����ד�F9��Y��G��u�&�9�!�'�m����M����\��T��*���
�l�m�n�w�}��������U��]�����h�}�'�6�9����HŹ��	��X�����
� �g�g��o�L���YӉ��P	��1��*��c�%�u�h��8�(���O����lU��1��U���&�9�!�%�f�;�(��M����l�N��*���1�
� �f�c��E��Yە��l��W�� ��b�
�g�:�w�0�(�������V��G�U���:�
�:�1��(�D��&���F��E1�����3�
�f�c�'�}�ϱ�&����9��h]�E���|�_�u�u�%�>��������9��R��]���
�8�`�
�2��G���ƿ�_9��G[�����a�e�|�_�w�}��������l ��V�*��i�u�7�8�%�8�ށ�����9����U���
�d�3�
�o�j����s���\��Q��*؊� �g�c�
�e�a�WǼ�����l��Q��G���%�u�;�u�:��A���&����l��d��Uʺ�0�3�:�
��(�E��&���F��E�����f�3�
�l�a�-�W���Y����
U��B1�C؊�g�n�u�u�8�8����&ǹ��lU��1��U��}�'�0�2��i����H�ӓ�F��SN����
� �f�a��o�L���YӉ��A ��@1��*��g�%�u�h��/����&����lT��1��U���u�8�
�`�1��G���	����F�G1�L���
� �l�d�'�}�J�������l��h�����
� �l�`�'�}�Ϭ�����l^��h�N���u�%�d�l�>�;�(��M����[�e��ۊ�9�
�0�:�����H˹��	��E�����f�a�%�|�]�}�W���Kù��l ��^�*��i�u�!�%�f�n����I�ѓ� F��<�����4�9�/�'�$�o����KĹ��]ǻN��*��
�
� �d�e��E��Yے��lW��h��D��
�f�:�u�6�:�F�������\��B1�Eڊ�g�n�u�u�'�l�E���&���� U��N�U¡�%�c�
� �n�l�����ƞ�]��h��*���:�
�
� �n�j����s���C9��1�����`�c�%�u�j�u����I����R��h�����;�0�
�;�����&����V��G\����u�
�
� �f�m�(��E��ƹF�N�����;�!�9�g���1���������R	�����b�c�e�u�w�l�^ϻ�
��ƹF�N�����;�!�9�g��f�W���	����ZW��B1�Aߊ�g�i�u�6�%�$�F���&����l��V ��'���0�
�9�
�9�.�B�������O��N����
�g�3�
�f�n����D�ί�A��1��*��c�%�u�;�w�<��������]��1��*��c�%�|�_�w�}�(�������T��h�I���6�'�,�3��o�D���Y����@��U�����d�d�%�|�]�}�W���&����W��N�U���u�u�u�4��2�����ޓ�u �������&�0�
�
�"�i�B���Q���A��N�����u�u�u�u�6�����&����lV��N����
�d�3�
�n�n����D�Ξ�]��h��*���&�f�'�2�c�j�W���Y����
T��B1�GҊ�g�n�u�u�'�i�(�������_��N�U�;�0�
�9��3��������W��N��ʡ�%�l�
� �d�m�(��B�����R����
�:�
� �e�l�(��E����^��V�� ��c�
�f�-�%�<�(���
����9��d��Uʥ��&�9�
��(�E��&���F��G1�� ����!��9�>�1�(��&����lT��1��]��1�"�!�u�c�f�W���	����F
��1��*��
�g�i�u�:�3�!�������9����U���
�g�
� �a�n����s���C9��D��*܊� �d�g�
�f�a�W���&����P9��T��]���<�0� �&�0�8�_���&����T��G]��@���n�u�u�%��.����&����S��N�U���
�:�<�
�2�)�Ǭ�
����F��P ��]���
�b�3�
�a��D��M����F�G1�����
�
�b�3��j�N���Y����K��z;�����
� �!�%�.�l�C�������_��F�U���;�:�`�|�]�}�W�������l��B1�Eފ�g�i�u�8�9�����I�ޓ� F��SN�����
� �d�l��o�L���YӖ��R
��^�� ��� �d�m�
�d�a�W���Y�����T�����d�
���w�5��������V9��^_�� ��`�
�g�e�w�}�F�������9F�N��U���4�g�d�
�"�l�Oׁ�J���F��a��*���3�
�d�g�'�}�J�ԜY���F��a��*ߊ� �
� �g�b��Dϩ�����V
��Z�*���g�e�
�g�g�}�W��PӃ��VFǻN��U���0�
�8�g��(�E��&����F�G1��؊�l�3�
�c�o�-�W��s���F�C��D���'�2�f�d�w�5��������CU��E��F���}�|�h�r�p�}����s���F�D�����c�3�
�c�g�-�L���YӖ��R
��1��*��e�%�u�h�]�}�W���Y����\��h��A��e�e�u�=�9�u��������9��P1�B���|�h�r�r�w�1��ԜY���F��a��*���'�2�f�c�l�}�WϮ�/����V��Z�����e�a�%�u�j�W�W���Y�ƭ�l��D�����b����w�5��������V9��^]�� ��l�
�g�e�w�}�F�������9F�N��U���4�g�`�
�"�o�Nׁ�K���F��a��*��
� �
� �d�d�(��E��ƹF�N�����;�!�9�f���1���?ӑ��]F��E�����
�a�3�
�f�h����P���A�R��U���u�u�u�%��1�(�������Q��UךU���
�4�g�g��(�(���K����CU�
NךU���u�u�%�6�9�)���&Ġ��u ��_��]���0�2�
�
�e�;�(��@����O�I�\ʰ�&�u�u�u�w�}��������l��h]�E�ߊu�u�
�4�e�o�(���J����CV�
N��*���&�
�#�`�n��_��T����\��XN�N���u�%��9��d����H�ޓ�F������g�
� �f�f��E��Y����G	�G�U���%��9�
��e����I�ԓ� F�d��U���u�4�
�:�$�����A����V��@��U �1�'�9�"�d�;�(��H����O�I�\ʰ�&�u�u�u�w�}��������l ��V�*��_�u�u�
�6�o�E���&����l��S��U���u�u�!�%�e����@Ĺ����YN�����
� �d�b��o�G���Y�����RNךU���u�u�
�
�"�l�Gށ�J���F��a��*���3�
�d�f�'�}�Jϭ�����Z��R�� �&�2�0�}��<�E��&����U��GZ��^ʠ�&�2�0�}�:��C���&����l��UךU���
�4�g�f�e����I¹��Z�=N��U���u�%�6�;�#�1�D݁�I����V��_��]���0�3�:�
��(�D��&���F�_��U���0�_�u�u�w�}�(���K����U��[����u�u�%��;��(���H����CT�
N�����2�6�#�6�8�u��������l0��1�����d�g�%�|�|�(�����θ�C9��h��D��
�d�|�_�w�}�(���K����U��]�����h�_�u�u�w�}�(���K����^��Q��F���%�u�=�;��3��������]	��E��F��}�|�h�r�p�}����s���F�G1��؊�
� �g�f��n�}���Y����_T��1��*���`�%�u�h�]�}�W���Y����V
��Q��@���%�u�=�;��/����K����S��h�E���u�d�|�0�$�}�W���Y����K��X
�����
�e�
�
�"�o�G߁�H���F��a��*ފ� �d�g�
�d�a�W���Y�����h\�����d�m�%�u�?�3�_���&����9��h_�G���}�|�h�r�p�}����s���F�D�����`�3�
�f�n�-�L���YӖ��R
��_�� ��l�
�g�i�w�)�(�������P�������1�%��9��m����M����M��Y�����!�%�l�
�"�o�Nہ�H����F�G1��؊�f�3�
�e�`�-�W��
����\��h����� �&�2�0������L����T9��W��^ʠ�&�2�0�}�:��C���&����l��UךU���
�4�g�`��(�D��&���FǻN��U���
�4�g�g�b�0����&����l��@��U �1�'�9�"�c�3����&����l��G��U��|�0�&�u�w�}�W���	����9��^�� ��e�
�f�_�w�}�(���K�ӓ�9��h\�@���u�h�_�u�w�}�W���*����U��X�����=�;�}�'�4�3�E���&����l��G��U��|�0�&�u�w�}�W�������_R��B1�Cڊ�f�_�u�u��<�E�������P��N�U���u�u�u�4��2�����ғ���YN�����
�0�
�b�f�m�W���H����_��=N��U���u�%�6�;�#�1�Eہ�I����l�N��#���
�
� �
�"�o�Bց�J���9F�N��U���6�;�!�9�e��1���?ӑ��]F��E�����
�
� �g�d��E��Y���O��[�����u�u�u�
�6�o�C�������]ǻN��*���g�c�3�
�a�k����Dӕ��l
��^�����'� �&�2�2�u�(���K�ߓ�V��\�U���;�<�;�1�#�-�B؁�����9��G�U���%��9�
��(�E��&���FǻN��U���-�
�:�0�#�/�(��&����lT��1��U���;�}�'�6�9����HŹ��V�
N��R���9�0�_�u�w�}�W���*����F9��^��F�ߊu�u�
�4�e�e����O�ӓ� F�d��U���u�;�"�0�a�;�(��N����D��F��*���1�
� �g�d��E��Y���O��[�����u�u�u�0��1�(���K����CU��N�����9�
�
� �b�n����D���F�N����c�3�
�c��l� ���Yے��lR��Q��Aߊ�g�e�u�u�f�t����Y���F���*���`�d�%�n�w�}��������_��B1�Fڊ�f�i�u�u�w�}�WϮ�/����V��Z�����e�a�%�u�?�3�_�������D9��Y�����e�m�%�}�~�`�P���Y����l�N��Uʥ��9�
�
�o�;�(��K����9F������&�3�
�m�o�-�W��s���F�V�����
�#�m�e� �8�WǪ�	����A��V�]���h�r�r�u�;�8�}���Y���R��X ��*���m�g�e�e�]�}�W���5����u	��{��*���!�3�
�`�g�-�W��
����\��h�����'�&�/�}�9�4����	����_��X�����&�3�
�`�e�-�^��P��ƹF��h�����:�
�:�%�$�;�(��K����[�N��U���4�
�:�&��+�F��������h_�*���f�l�
�f�g�}�W��PӃ��VFǻN��U���8�
�`�
�"�n�@ށ�H���F��Y��ۊ� �g�`�
�e�a�WǺ�����l��X��*���g�g�
�f�/�/��������_��G�U���%�;�!�<��(�D��&���F��R�����0�:�
�
�"�n�Nف�JӞ����T�����d�d�n�u�w�-��������T��h�I���1�9�!�1�-�/�������� W��N��ʴ�
�:�&�
�!��^�ԜY�Ƽ�\��Q��@ߊ�g�i�u�!��2����������Y�����:�&�
�#��h�W���������h_�*���c�d�%�|�l�}�WϮ�����lW��1��U��&�1�9�2�4�+����Q����V��G1�����9�c�f�|�z�.����Q���� R��B1�B܊�d�|�_�u�w��(���K����CU�
NךU���u�u�%�6�9�)����Hӑ��]F��Z��D���2�f�l�}�~�`�P���Y����l�N��Uʴ�
�:�&�
�!��L���Y�����1�����
� �b�f�'�}�Jϭ�����Z��R��§�&�/�}�<�9�9����&¹��lQ��h�Y��|�_�u�u�'�.�(ށ�����l��S�����:�<�
�0�#�/��������R��X ��*���g�g�u�u�9�4����?����U��W��G���_�u�u�u�w�2�F���
����lW��1��U��&�1�9�2�4�+����Q����I��^	��¥�&�
� �d�b��E��K����9F���D���
�f�a�%�w�`��������l��C�� ���2�0�}�%�4�3����H����M��Y������
�0�
�`�d�^�ԜY���F��D\��*���!�3�
�e��l�K�������T��A�����0�<�0�&�0�8�_���K�ד�F9�� 1��\��|�n�_�u�w�2�E�������9��R�����9�2�6�#�4�2�_���������T�����d�
�|�~�"�.����Q�ԓ�l ��W�����n�u�u�u�w�-�݁�����F9��V��D��u�!�
�:�>�����۔��Z��D�����:�g�3�
�d�n����J���9l�N��؊� �d�c�
�e�a�W���&����P9��T��]���<�;�1�4��2�����ԓ�F�B �����}�g�'�2�d�j�^��Y����Q9��Q��Gߊ�f�i�u�u�w�}�WϷ�����l ��]�����=�;�}�8��m����I¹��V�
N��R���9�0�_�u�w�}�W���&����U��Y��F�ߊu�u�7�4�$�:�(ށ�����9��R��]���
�
� �d�d��EϿ�ӗ��U��[�����_�u�u�7�6�.����&����U��G\��H���
�
�d�'�0�n�C����ƽ�lW��R	��M��n�u�u�$��.����L����W��h�I���'�<�<�
�"�o�@؁�KӇ����C1��*��b�%�|�_�w�}����
����9��h\�L���u�h�}�
��n����A�ғ�F��SN�����
�0�
�e�f�f�W�������@��hW�� ��a�
�g�i�w�/����&����R��G\�����7�!�g�'�0�i�G���s���B��B1�@ي�f�i�u�u�w�}�WϷ�����V�� [����u�!�%�d��(�F��&���F�_��U���0�_�u�u�w�}����A����W��h����u�7�!�3��l�@���Y����l0��1�*���f�d�
�g�n�9� ���Y����F�E1�����l�
�g�i�w�)���&���� U��N��ʡ�%�`�
� �a�h����s���A9��Q��D���%�u�h�w�u�*�������� Q��B1�@ފ�d�h�4�
�8�.�(���&����_��_�����u�
�
� �e�j�(��E���F��R �����d�`�'�2�c�h�W���	����@��A\��E���9�0�w�w�]�}�W���&����U��G\��H���w�"�0�u�#�-�F�������V��
N��*���&�
�#�d�g�}����[����F�E1��D���
�m�
�g�k�}��������E��X�����
�<�=�}�9�4��������]��[�*ٓ�������[�������V��Y�����r�r�s�!�'�k�(���A�ߓ�N��_�����:�e�|�|�l�}�WϬ�/�ғ�F9��_��G��u�!�
�:�>�����ە��]��C��Mފ� �g�`�
�f�}�W�������^��1��*��f�%�|�n�w�}����L����P��h�I���!�
�:�<��8����
����WN��G1�*���g�b�
�d�w�}����ے��l^��Q��C���%�|�n�u�w�/�!���&����l��S�����:�<�
�0�#�/��������[��Y�����4�
�:�&��+�C���?����u ��q(��Y���<�!�2�'�"�.����Q���F��G1�*���d�`�
�d�d�p�W������O�UךU���
� �d�d��o�K�������9��h_�E���u�;�u�8��e����K�֓�O��N�����<�
� �b�n�-�W��Q����T��Q��Eߊ�d�:�u�
��(�A���	����F�E1��؊� �g�b�
�e�a�WǪ�	����l ��_�*��:�u�
�
�"�o�B؁�K��ƹF��h��F���
�m�a�%�w�`�_���&����A��^�U���'�f�3�
�o�d����s���A9��^Z�� ��a�
�g�i�w�)���M����lR��N��U���
� �f�f��o�L���YӔ��l��B1�Fފ�g�i�u�!�'�k�(���H����CW��EN�����g�c�%�|�]�}�W���H����R��h�I���!�%�d�m�1��C���	�ƴ�AF��h�����#�
�|�_�w�}��������9��R��]���
�f�
� �o�n�����ƭ�l��D��ۊ�|�_�u�u�2�n����O¹��Z���*��
� �m�f�'�}����	����@��A_��\�ߊu�u�0�b�1��C���	���N��X��2��� �
�'�4�2���������l ��]�*��-�'�4�
�8�.�(���&����F�E��*���f�a�
�g�k�}����H�ѓ�V��Z����4�
�:�&��+�(���s���A��h��F��
�g�i�u�#�-�F�������V��N��ʴ�
�:�&�
�!��^�ԜY�ƾ�E9��h_�A���u�h�}�8��o����J�Г� F��EN��*���&�
�#�
�~�W�W�������CW��Q��C���%�u�h�w�u�*��������l ��h"�����'�2�f�e�j�<�(���
����9�������w�_�u�u�2����&����^��G\��H���0�
�8�`�1��E���	�ƭ�WF��G1�*���d�g�
�f�l�}�Wϭ�����T��Y�����b�`�%�u�j�u��������U��[�����:�u�%�6�9�)����H��ƹF��R����
� �d�m��n�K���Y���F��h8��G���3�
�g�e�'�}����Q����G��1��*��f�%�}�|�j�z�P������F�N�����!�%�
� �f�k�(��s���@��C��F���
�g�b�%�w�`�_���&�ד�F9��\��Fʭ�'�4�
�:�$��ށ�P���F��[1�����3�
�f�f�'�}�J�������CS��B1�BҊ�g�4�1�&�;�)��������
Q��G�U���&�9�!�%�b���������F9��V��G��u�!�%�f��8�(��HӉ��Z��1����c�|�_�u�w�8�(���Hƹ��lW��1��U��_�u�u�u�w�����J����T��h����u�&�9�!�'�i����J�Փ�N��S��D���0�&�u�u�w�}�Wϭ�����T��B1�Mӊ�f�_�u�u�2����&���� W��G\��H���w�"�0�u�$�:����K����lU��G��U���;�1�4�
�8�.�(���K����F��D��E��u�u�&�9�#�-�@ځ�����R��B1�Aӊ�g�i�u�<�:�n����M�ѓ�F����B���
�a�f�%�~�W�W�������CW��Q��F���%�u�h�}�2����&���� W��G\�����8�
�
� �f�e�(��B�����h��D���1�8�'�4��(�E��&���F��R����`�1�8�'�6����Mʹ��	��C��Bӊ� �g�d�
�e�f�W���
����^��h��D��
�g�i�u�#�-�O݁�����9�������g�
�:�
�"�l�D߁�K��ƹF��R����
� �d�a��o�K�������9��h_�G���u�;�u�0��0�Fׁ�����9��UךU���0�
�8�d�1��B���	���l�N��Uʥ�<�
�!��%���������F9��^��Dʢ�0�u�&�9�#�-����L�ד�N��S��D���0�&�u�u�w�}�WϷ�&����\��h�����:�
�:�%�$�;�(��M����9F���*���g�
� �d�c��D��Y���F�<�����4�9�:�0�����Kù����YN�����8�d�
� �f�i�(��I���W����ߊu�u�u�u�2����@ǹ��l�N�����%�d�3�
�b�i����D���F�N�����
�9�
�0�8����Iù����YN�����8�d�
� �f�i�(��I���W����ߊu�u�u�u��l�(�������9��d��Uʦ�9�!�%�g�1��N���	���N��G1�*���
�l�m�-�%�<�(���
����9��d��Uʦ�9�!�%�f�1��N���	���N��GZ�� ��c�
�g�4�3�4��������S��d��Uʦ�9�!�%�a�1��N���	���N��G1�*���
�l�m�4�3�4��������S��d��Uʦ�9�!�%�`�1��G���	���l�N��Uʥ��9�
�
�"�o�Aف�Jӑ��]F��Z��G���
�e�f�%��t�J���^�Ʃ�@�N��U���%��9�
��8�(��A���F��[1����
�0�:�2�9�;�(��K����[�C��Lӊ� �f�`�
�e�2�W���&����U��[�����_�u�u�0��0�Eف�����
9��R�����u�u�u�0��0�Eځ�����9�������0�
�8�l��8��������V��h�E���u�d�|�0�$�}�W���Y����l0��1�����f�l�n�u�w�.����	����W��E	��*���f�e�
�g�k�}�������� 9��Z����� �f�m�
�e�2�W���&����U��X�����_�u�u�0��0�E؁�����9��R��]���
�
�0�
�`�l��������]��[��D��u�u�&�9�#�-�O���&����l��S�����
� �g�e��o��������A��Y�\�ߊu�u�0�
�:�o�(���N�ӓ� F�d��U���u�!�%�d�b�;�(��&����[����*���3�
�f�
�e�m�W���H����_��=N��U���u�%�6�;�#�1�Fׁ�B�����h��G���
�`�a�%�w�`�_���&����U��Y�����:�u�%�6�9�)����H��ƹF��R����
� �b�f�'�}�J�������l ��]�����:�u�%�6�9�)����H��ƹF��R����
� �b�l�'�}�J���,����}%��h��@���%�u�;�u�2����&����U��G�U���&�9�!�%�e�;�(��@����[�D�����d�'�2�f�b�}��������9��P1�F���_�u�u�0��0�D܁����� 9��R�����u�u�u�
�6�o�A���&����l��@��U¦�9�!�%�g�1��A���	����[�I�����u�u�u�u�w�.����	�ߓ�V��Z����u�0�
�8�d����Nù��Z���*��
�0�
�m�c�%�Ͽ�&����G9��1�N���u�&�9�!�'�h����O�ӓ�F�F�����%�d�'�2�d�h�W���Y����G��1��*��e�%�|�_�w�}��������U��V�����h�_�u�u�w�}�(���K�Г�F9��X��Gʢ�0�u�&�9�#�-�B���&����l��G��U��|�0�&�u�w�}�W���
����^��h��D��
�f�_�u�w�8�(���JĹ��lQ��h�I���<�8�d�3��i�(������^��1��*���
�g�n�u�w�.����	�ޓ�F9��1��U��}�8�
�f��(�O���	�ƣ���hX�����3�
�`�
�e�f�W���
����^��h��L���%�u�h�}�:��O���&����CT��Y
�����8�f�
� �n�n����s���@��C��*���f�a�
�g�k�}����&����W����U���
�8�g�3��h�C���P���F��[1�����3�
�b�
�d�a�W���Y���4��P�����:�0�
�
�"�e�@���Y����N��[1�����3�
�c�
�e�m�W���H����_��=N��U���u�0�g�3��o�(��s���@��C��D���
�l�
�f�k�}�W���Y����R��1�����'�&�g�3��o�(��������h��Fӊ� �l�l�%��t�J���^�Ʃ�@�N��U���%�d�l�<��(�N���	��ƹF��R����
� �d�b��o�K�������
9��P1�C���:�u�%�6�9�)����H��ƹF��R����
� �d�l��o�K�������l ��Y�*��4�1�<�;�0�l����J����l�N�����%�a�3�
�`�e����D�θ�C9��h��*��l�4�1�<�9�:�F�������O��N�����!�%�`�3��d�G���Y���F�N�����9�
�
� �f�e�(��������hY�����m�`�%�}�~�`�P���Y����l�N��Uʥ��9�
�l�1��A���	��ƹF��R����
� �d�d��n�K���Y���F��R����
� �d�e��n� ���Yە��l��[�����'�4�
� �f�m�(��I���W����ߊu�u�u�u��<�E��&����^��G]�U���&�9�!�%�`�;�(��I����[�C��FҊ�0�
�m�d�/�/��������_��G�U���&�9�!�%�o�;�(��H����[�C��G���
�l�`�%�w�3�W���	����T9��]����u�0�
�8�c����JĹ��Z���ي� �g�e�
�e�%�Ͽ�&����G9��1�N���u�&�9�!�'����Mƹ��Z�=N��U���u�;��'�8��W����ο�_9��G]�� ��a�
�g�e�w�}�F�������9F�N��U���
�8�d�3��h�A���B�����h��@ڊ� �g�a�
�e�a�WǬ�Ĺ��lT��1��U���u�0�
�8�c����JĹ��]ǻN�����8�`�
� �e�k�(��E����\	��O)��:����0�!�'������&����lT��1��U���u�6�%�b�9�)����M�ӓ�O��N�����!�%�g�3��i�@���Y���G�� W�� ��d�
�g�4�3�.����	�ד�F9��_��G��u�u�&�9�#�-�D���&����l��S�����!�%�m�
�2�2��������U��N��ʴ�
�:�&�
�!��^�ԜY�ƿ�_9��G[�����a�`�%�u�j�u����I����R��h����&�9�!�%�d�;�(��@����l�N�����%�a�;�!�1��B���	���N��[1�����3�
�g�f�'�}����	����@��A_��\�ߊu�u�0�
�:�h�(���K����CU�
NךU���u�u�%�6�9�)����Kӑ��]F��R�����
�0�
�e�g�m�W���H����_��=N��U���u�%�6�;�#�1�D��s���@��C��C���
�c�e�%�w�`�}���Y���@��C��@���
�c�f�%�w�5��������WW��B1�G݊�g�e�u�u�f�t����Y���F���*���g�e�
�f�]�}�W���&����9��h\�M���u�h�_�u�w�}�W�������l
��h]�����}�0�
�8�b�����I���F�_��U���0�_�u�u�w�}��������EU��d��Uʦ�9�!�%�m�1��E���	���N��G1�*���f�`�
�g�/�/��������_��G�U���&�9�!�%�n�;�(��O����[�C��D���3�
�g�`�'�}��������CS��Q��G���%�|�_�u�w�8�(���L����T��h�I�����
���8�(��KӇ����h��L���
�g�g�%�~�W�W�������CP��Q��G���%�u�h�}�2����J����\��Y1��*��g�%�u�:�w�-��������lW�=N��U���
�8�c�
�"�n�Nہ�K�����h_�*���f�c�
�g�6�9��������l ��\�*��n�u�u�&�;�)��������P��N�U¦�9�!�%�b��8�������� U��h����4�
�:�&��+�(���s���@��C��F���
�f�g�%�w�`�_���&����U��X�����;�u�0�
�:�k�(���J����CT�=N��U���
�8�c�3��h�E���Y���G��[�����a�a�u�;�w�8�N���&����l��d��Uʦ�9�!�%�
�"�l�Aہ�J���9F�N��U���
�l�3�
�g�l�������G��1��*��c�%�}�|�j�z�P������F�N�����:�&�
�#�c�m�}���Y����G��h��F��
�g�i�u�f�}����Q����Z9��E1�����
�0�
�d�w�}��������ET��N�����e�n�u�u�$�1����J����\��Y1��*��`�%�u�h��0�(؁�����W��EN�����0�
�b�m�l�}�Wϭ�����
9��h_�G���u�h�}�8�����OŹ���������!�9�d�d�l�}�Wϭ�����l ��[�*��i�u�!�%�f�n����M�ӓ�F��SN��Ҋ�0�
�d�f�l�}�W���Yӕ��R��1����� �`�d�%�w�`��������l��C�����/�}�<�;�3�.�(���&¹��lS��h�Y��|�_�u�u�$�����&����U��N�U���u�u�u�!�'�n�(���L�ד�F��R ��$���
��
�
�"�h�B���Q���A��N�����u�u�u�u�#�-�C߁�����l��=N��U���u�=�4�!�4�.�(���H����CW�
N�����2�6�#�6�8�u����ە��]��D����� �d�`�
�d�q�E���s�����V�����e�`�%�u�j�W�W���Y�Ƹ�C9��Q��E���%�u�=�;���9���:����lU��F�U���d�|�0�&�w�}�W���YӒ��lW��B1�@ڊ�g�_�u�u�>�3��������U��^�����h�_�u�u�w�}����@����Q��h����u�&�9�!�'�i����N�ޓ�N��S��D���0�&�u�u�w�}�Wϭ�����U��B1�Lي�g�_�u�u�>�3��������]	��Q��M���%�u�h�}�>�3��������U��^�����:�u�%�6�9�)����H��ƹF��^	�����2�
� �d�o��D��Y���F���*���3�
�l�f�'�}����Q����G��1��*��l�%�}�|�j�z�P������F�N�����!�%�f�3��d�C���B�����Y1�����
�:�
� �e�i�(��E����Z��V����� �d�m�
�d�%�Ͽ�&����G9��1�N���u�&�2�7�#�;�(��H����[��h8��G��
� �f�d��o�D�������U��d��Uʡ�%�e�3�
�`�j����D�΢�D��Y��*ۊ� �d�d�
�d�<�ϭ�����T��B1�B܊�g�n�u�u�#�-�F���&����l��S�����3�:�
�
�"�l�D݁�KӉ��@��h�����d�;�!�3��e�E���P���F��G_�����l�`�%�u�j�u�����ד�F9�� Z��Gʴ�1�&�9�!�'�j����@�֓�O��N�����f�3�
�g�b�-�W��Q����Z��^��*���g�l�
�f�8�}����O����T��h�N���u�!�%�a�1��N���	���N��G]�*���:�2�;�3��d�N���Y����R��X ��*���
�|�_�u�w�0�Fځ�����9��R��]���0�2�a�
�2�2����¹��lT��1��U���!�%�l�
�"�o�A݁�K��ƹF��Z�*���f�c�
�g�k�}����K����^	��V �� ��`�
�g�-�%�<�(���
����9��d��Uʡ�%�b�3�
�f�l����D�ή�^��RZ�����'�4�
�g�1��F���	�ƣ���hW�����d�d�%�|�]�}�W���H˹��lU�� 1��U��&�1�9�2�4�+����Q����T����%���:�
�|�~�"�.����Q����_T��1����`�|�n�u�w�)�ށ�����9��R��]���f�`�1�8�%�<�(���H����CT��X�����;�!�9�d�f�f�W�������U��_�����h�}��3��i�G���Y����A��Q��F���%�|�_�u�w�0�D�������T��Q��F���%�u�h�}�:��A���&����l��X�����8�d�
� �f�o�(��B�����^�����
�4�!�3��d�(��E��ƹF�N�����;�!�9�d��}����Q����l/��h��F���%�}�|�h�p�z�W������F�N��*���&�
�#�g�f�W�W�������l��X�����
�c�a�%�w�`�_���&����U��[�����'�&�9�!�'�j����J����l�N����
�4�!�6�$����N����[�N��U���4�
�:�&��+�E������7��y1��6���3�
�e�
�e�m�W���H����_��=N��U���u�%�6�;�#�1�F݁�B�����_�����'�4�
� �e�j�(��E����lU��^1��*��f�%�u�'�5�0����I����\��Y1�����g�b�%�|�]�}�W���J�ד�V��P�����l�l�%�u�j�u�(���¹��lT��1��U���7�8�'�0�g�9��������l ��W�*��n�u�u�!�'�o�(�������l ��_�*��i�u�%�f��o����H�Փ�F�������a�
�0�:�0�3�݁�����9��UךU���8�f�3�
�b�k����D�ο�_9��G_�����f�g�%�u�%�.����	�ғ�\��B1�Mڊ�g�n�u�u�#�-�(���H����CT�
N�����2�7�!�'�0�n�F����ƿ�_9��G\�����l�l�%�|�]�}�W���L����V��h�I���:�0�3�:��(�E��&����AF��P �����;�;�!�3��m�F���P���F��GX�� ��e�
�g�i�w�?��������V��h����&�9�!�%�`�;�(��O����l�N��݊� �d�l�
�e�a�WǪ�	����W��E	��*���d�l�
�g�/�/��������_��G�U���!�%�
� �o�l����D�Π�lW��B1�B���u�;�u�0�e�;�(��&���9F���L���
�b�d�%�w�`�_���&����9��P1�@���'�&�9�!�'�o�(���&����T��G\����u�8�
�e��(�D��&���F�N����� �
�&��$���������R��E��A��u�u�%�6�9�)����K�Ʃ�@�L�U���!�%�d�d�1��E���	���D��������6�
�4�2���������^��R	��E��h�4�
�:�$��܁�PӃ��VF�UךU���8�
�e�
�"�n�Aځ�K���W�@��U �
�&��&��)��������9��P1�F���u�%�6�;�#�1�D��Y����D��d��Uʡ�%�d�f�3��i�B���Y���D��_��]���;�1�<�
�#���������9��h]�G���|�i�&�2�2�u��������O�R��U��n�u�u�!�'�l�C���&����l��S��9��� �,� �
�g����Oƹ��U��S�����|�_�u�u�:��Gׁ�����9��R�����
� �d�c��o�F�������W��d��Uʡ�%�d�l�3��k�A���Y����\��Q��F���%�}�d�1� �)�W��B���F���*���3�
�d�m�'�}�Jϭ�����Z��R��§�&�/�}�<�9�9����Hʹ��lW��1��\��|�n�_�u�w�0�(��&���� W��N�U���2��d�3��o�(��O���F��@ ��U���_�u�u�8��l�(���M�Փ�F������d�3�
�g��l�B���Y�ƨ�D��^����u�8�
�d��(�B���	�����h8��*���a�`�%�}�o�p�FϺ�����O��N�����d�c�3�
�a��F��Y����P��B1�D���}�m�x�d�3�*����P���F��G1�B���
�m�
�d�k�}����@����^��G\��M���d�1�"�!�w�t�}���Y����W��Q��D݊�f�i�u�4���(���M�ӓ� N��h�����}�;�<�;�3�)���&����l ��_�����u�:�;�:�#������ι�@��R
�����c�6�&�
�"�k�D���P����[�������2�'� �&�0�8�_���&�Г�R��Q��Dي�d�|�h�e�6�9��������AN��D�����8�
�c�6�$����J����Z�G�����w�w�_�u�w�0�(��&����W��N�U���
�a�3�
�d��E��T����\��XN�N���u�!�%�d��(�F��&���F��S1�����#�6�:�}�?�;�(���ۓ��Z��SF����
� �d�e��l�[�������V��Y�����r�r�s�&��0�(�������V��h�F���u�:�;�:�g�t�^��Y����^��^�� ��d�%�u�h�]�}�W���Y����\��h��*���=�;�}�8��h����Mƹ��V�
N��R���9�0�_�u�w�}�W���	¹��lP��h����u�8�
�g��(�A���	�����h�����0�!�'�'�$�'�_���������h_�*���c�d�%�|�b�t�L���YӒ��lW��h��C���%�u�h�&�3�1��������AN��^�����!� �&�2�2�u��������ES��(��3������|�#������ι�@��R
��E���u�8�
�g��(�A���	����W��X����|�|�n�u�w�)���L����V��G_��Hʥ��9�
�
�"�h�D���Q���F��@ ��U���_�u�u�8��o�(���H����CU�
N��#���
�
� �d�c��E��Y����G	� G�U���!�%�d�b�1��Dځ�M���uT��h��A���%�}�d�1� �)�W���s���G��\�����b�
�a�i�w�0�(�������9��_����!�u�|�_�w�}����K����W��h�I���d�u�=�;��4��������l ��^�*��u�u�<�;�3�<�(���
����T��G�����u�e�n�u�w�)���I����W��G]��Hʥ�&�
�
� �`�j����Hӂ��]��_����u�8�
�f��(�O���	�����1�����l�
�g�d�w�2����H����F�C��D���3�
�e�b�'�}�JϮ�
¹��U��Y��G��u�:�;�:�f�t�}���Y����U��Q��D���%�u�h�%��1�(�������^��F�X��1�"�!�u�~�W�W�������9��h\�F���u�h�%��;��@���&����l��]�����:�f�|�_�w�}����Jʹ��lT��1��U��%��9�
�`�;�(��A����V��X����|�_�u�u�:��D���&����CW�
N�����
� �f�l�'�u�E��Hӂ��]��G�U���!�%�d�d�1��D���	�����V��Aۊ� �g�f�
�d�o�W������ O��N�����d�g�3�
�d�d����D�ή�\
��p+�� ���'�4�0�
�%�����
����U��h�Sʷ�:�
��e�"���������l#��V��*���g�`�
�g�l�}�WϪ�	����l ��Y�*��i�u�-�
������&����Z��h_�*��� �g�m�
�e�o�W���Y����G	�UךU���8�
�a�3��l�A���Y����G��X	��*���!�'�&�2�2�u��������EW��q+�U���<�;�1���8�(��@����F�C��D���3�
�m�f�'�}�Jϸ�	����2��B�� ���%�,�d�b��;�(��@����W�_�����:�e�n�u�w�)���A���� R��h�I����9�
�:��2���H���� R��h�F���u�u�:�;�8�m�L���YӒ��lW��h��F��
�f�i�u��1�(���&����lT��h��F��
�`�f�u�8�3���P���F��G1�*���d�c�
�g�k�}�F������@��R
��G���2�f�b�|�i�.����Q����\��h��G��|�u�9�0�u��}���Y����P��Q��A���%�u�h�<��)�1���5����V��Q��A���%�}�d�1� �)�W��B�����h_�����d�`�%�u�j�.��������V��EF�����}�%�6�;�#�1�F݁�<�����Y��3؊�0�
�b�l�~�W�W�������l ��_�*��i�u�d�u�?�3�_�������^��1��*��`�%�|�k�$�:����	����@��A_��F���u�9�0�w�u�W�W���Y�Ƹ�C9��h�����
�d�d�%�w�`��������l��C�����/�}�<�;�3�)���&����U��G\��F���n�_�u�u�:��O���&����l��S��E���=�;�}�
�2�(��������R��N�����:�&�
�#�c�m�W�������l�N����
� �d�b��l�K�������U��]�����a�x�d�1� �)�W���s���G��1��*��e�%�u�h�$�9��������G	��B �����}�%�6�;�#�1�F݁�O���F��P ��]���'�2�f�b�~�f�W�������9��h_�C���u�h�&�1�;�:��������A��M�����;�1�$�
�$�4��������V��G�A���_�u�u�8��l����Iƹ��Z�D�����6�#�6�:��3����ے�� V��T��*���!�3�
�l��n�W�������V��O��*���f�l�%�|�l�}�WϪ�	����U��V�����h�w�w�"�2�}�����μ�@W��B1�@ފ�g�u�u�<�9�9��������_��h]�\ʰ�&�u�e�n�w�}����K����lW�� 1��U��!�%�l�3��m�F���Q���W��X����n�u�u�!�'�o�(���H����CW�
N�����2�6�#�6�8�u����ۓ��Z��SF��ۊ�4�!�3�
�d�d����L���9F���*���3�
�d�m�'�}�JϪ�	����U��_�����a�x�d�1� �)�W���s���G��X�� ��e�
�g�i�w�)�(�������P�������<�=�}�<�9�9����/����V��h�Y���<�!�2�'�"�.����Q���F��G1�*���d�e�
�d�d�p�W������O�UךU���8�
�b�3��i�G���Y���D��_��]���;�1�%�&��(�F��&���F��P ��]���6�;�!�9�f��A�������V�=N��U���
�m�3�
�f�h����DӋ��l0��B1�FҊ�f�!�
�;�2�8�_���������h_�����
� �d�a��l�^Ϻ�����G	��Y�����;�<�;�1�#�-�Fׁ�����F9��_��D���u�=�;�}�8�4����ۓ��Z��SF����
�4�!�3��l�F���P���F��SN��*���0�0�}�;�>�3�Ǫ�	����P��h��D��
�d�|�h�d�}����[����F�C��Gӊ� �d�`�
�f�a�W���&����P9��T��]���<�0� �&�0�8�_���K����G9��h_�M���|�`�|�n�w�}����Kʹ��G9��h_�E���u�h�}�8��j����M�֓�F��EN��*���&�
�#�
�~�W�W�������U��[��D��u�!�
�:�>�����۔��Z��B �����}�-�
�8�����L����W��UךU���8�
�e�3��i�C���Y���D��_��]���2�g��d�1��C���	���R��X ��*���a�e�u�9�2��U�ԜY�Ƹ�C9��h��D��
�g�i�u�f�}����Q����l ��]�*��h�4�
�:�$�����J����_��^�����u�8�
�g�1��G���	���N��G1�����f�b�u�'�"�9��������V��h�N���u�!�%�f��(�F��&���F��V ��D���9�:�0�
���C���&����l��O�����:�&�
�#��t�}���Y���� R��B1�B܊�d�i�u�8��k����H�ӓ�N��N����!�u�|�_�w�}����L����V��h�I���<�;�2�'�0�n�B����ƭ�l��D��ۊ�|�_�u�u�:��A���&����CW�
N�����2�6�#�6�8�u����ۓ��Z��SF�����%��d�3��i�(��U���l�N����
� �a�b�'�}�J���	����@��A_��U���8�
�d�
�"�i�D���P���F��G1�*���a�f�%�u�j��Uϩ�����^��\�� ��d�%�u�u�'�>��������O��[��W���_�u�u�8��d����H¹��Z�D�����6�#�6�:��4��������]��[�*���|�~�&�2�2�u�E�������
9��G�U���!�%�f�3��m�A���Y���D��_��]���'�2�f�b�w�}��������EW��X�����u�e�n�u�w�)���&����Q��N�U���
�:�<�
�2�)�ǫ�
����WN��h�����#�g�d�|�z�(�����Ί�lW��B1�L���|�n�u�u�#�-�Cށ�����l��S��D���=�;�}�g�f�;�(��&�����T�����d�
�e�u�;�8�U���s���G��\�� ���`�%�u�h�u�� ���Yۓ��Z��SF��*���
�
� �`�d�-�^������]��V�����
�#�g�f�~�}����[����F�C��Aي� �d�m�
�d�a�W���Y�����T�����c�e�"�0�w�)���&����Q��G\��\��r�r�u�9�2�W�W���Y�Ƽ�\��B1�Mڊ�g�_�u�u�:��C���&����CT�
N��Wʢ�0�u� �&�0�8�_�������l ��\�����i� �&�2�2�u��������EW��\��U���0�w�w�_�w�}����L����S��G_��Hʦ�1�9�2�6�!�>����������^	��¦�
�8�
�
�6�)����J¹��J��G�U���!�%�a�
�"�h�F���Y����G��X	��*���!�'�&�<�#�/����
����WN��Y1��C���
�m�
�f�{�2��������]��Y��R��s�!�%�a��(�B���	����W��X����|�|�n�u�w�}�WϪ�	����U�� W��D��u�!�
�:�>�����۔��Z��D�����8�
�d�
�"�h�F���P����]ǑN�����a�
� �d�n��F��Y����_	��T1�����}�0�<�0�"�.����Q����U��B1�M܊�f�y�a�|�]�}�W���&�ߓ�F9��1��U��&�1�9�2�4�+����Q����G9��Q�����;�1�!�%�c����@������^ ����� �&�2�0��m�W�������lW��V�����f�
�d�f�z�}�������O�=N��U���
�
� �f�d�-�W������e9��h]�*��c�u�u�u�8�3���B�����h[�����e�
�g�i�w�l�W����ο�T����*���3�
�d�
�e�}�W�������C9��Y����
�c�|�0�$�}�G��Y����^��1��*��m�%�u�h�$�9��������G	��D�����2�!� �&�0�8�_�������l
��1��3�������~�)�(�������F��P ��]��u�u�8�
�o�;�(��M���� W�
�����e�|�|�n�w�}����L����lP��h�I���!�
�:�<��8����
����WN��h�����#�g���w�}����۠��9��hZ�*��|�_�u�u�:��D���&����CT�
N��Wʢ�0�u�&�2�2�u�E�������
9��N����0�}�%�6�9�)���&�����RN��W�ߊu�u�8�
�c�;�(��&���F��S1�����#�6�:�}�>�3�ǿ�&����G9��\��0���~�&�2�0��o�F���&����CT�d��Uʡ�%�`�
� �a�h����D������YN�����1�!�%�`��(�A���	�����Y�����:�&�
�#�e�n�^������D��N�����`�
� �c�b�-�W��[����[�������!�g�3�
�`��E������]��[�*���0�&�u�d�l�}�WϪ�	����U��Z�����h�&�1�9�0�>�����ξ�@�������1�$�
�&�>�3�D���&����l��_�\�ߊu�u�8�
�o�;�(��&���F��S1�����#�6�:�}�9�4�������� 9��D�����3�
�`�
�d�}�W���������h8��*���a�b�%�|�l�}�WϪ�	����U��Y��G��u�d�u�=�9�u����ۖ��9��Q��M݊�g�u�u�<�9�9��������_��h]�\ʰ�&�u�e�n�w�}����L����V��h�I���d�u�=�;��3����ە��R��Q��E���%�|�i� �$�:����	����@��A_��F���u�9�0�w�u�W�W�������l ��\�����h�&�1�9�0�>�����ξ�@�������1�%�&�
��<����&����CW�Z��N���u�!�%�c��(�F��&���F��a��*؊� �d�g�
�d�o�W������ O��N�����c�
� �m�f�-�W��
����\��h�����&�<�!�'�0�)�����Ρ�]9��1��*��
�f�y�:�>�)��������]��^��Sʡ�%�c�
� �o�j����H����\��XN�\���n�u�u�!�'�k�(���H����CW�
N��#���
�
� �d�e��D��T����\��XN�N���u�!�%�c��(�O���	���D�������<�;�1�%�$��(���N�ѓ�O������4�
�:�&��+�E��P�Ʃ�@�L�U���!�%�c�
�"�e�N���Y����G��X	��*���!�'�'�&�-�u��������\��1����� �m�f�%�~�h�^��Y���F��Z��C���&�
� �c�d�-�W��
����\��h�����'�&�/�}�>�3�Ǫ�	����U��Y��G���g�|�_�u�w�)���&����S��G]��Hʥ��9�
�
�"�l�B߁�K����W	��C��F��u�u�!�%�a����H����[�L�����}�4�2�g��n����A����[��G1�����9�`�
�|�2�.�W��B�����hX�����3�
�`�
�e�a�WǪ�	����U��Y��Gʭ�'�4�
�:�$��ށ�P���F��G1�*���l�l�%�u�j��Uϩ�����\��1��*��
�g�h�4��2�����ԓ�O��[��W���_�u�u�8��d����N�֓�F�F�����
�9�
�;�$�o�ށ�L����Q��h����4�
�:�&��+�(���s���G��1��*��d�%�u�h�u�� ���Yۓ��Z��SF��*���
� �d�`��n�W�������V��G1�����9�d�
�m�~�8����I��ƹF��Z��E���
�m�`�%�w�`�_���&�ޓ�V��_����;�0�3�:�����Lù��]ǻN�����d�3�
�m�`�-�W��Q����T9��E��F��u�:�u�%�4�3����H���9F���*���3�
�d�
�c�a�W���&�ד�F9��1��]��1�"�!�u�~�W�W�������l ��]�*��i�u�d�u�?�3�_�������l0��1�*���
�l�c�u�w�4��������]��[�*���u�9�0�w�u�W�W�������l ��_�*��i�u�!�
�8�4�(�������V��RF�����0�}�7�4�$�:�(ځ����� 9��B�\��u�u�!�%�`����IĹ��Z� �����7�!�g�3��l�N���Y����R��X ��*���
�|�_�u�w�0�(������� Q��N�U¦�2�7�!�3��l�F���Y����R��X ��*���
�|�_�u�w�0�(�������Q��N�U��u�=�;�}�>�3�Ǯ�/����W��B1�F܊�f�u�u�<�9�9��������_��h^��U���0�w�w�_�w�}����A����U��h�I���}�:�9�-����������l)��r�����3�
�f�f�'�}�W�������)��h)�����
�'�� �;�l����J�ד�O��������!��2�)����&����_9��Q��G���%�|�_�u�w�0�(�������_��N�U��u�=�;�}�:��O���&����l��
N��*���&�
�#�
�~�8����I��ƹF��Z��*���f�l�%�u�j��Uϩ�����^��h��F���%�u�u�%�4�3����O������RN��W�ߊu�u�8�
�g�;�(��L����[�L�����}�8�
�m�1��D���	���R��X ��*���
�|�0�&�w�m�L���YӒ��l^��Q��A���%�u�h�w�u�*��������9��h\�L���u�u�%�6�9�)����N�Ʃ�@�L�U���!�%�m�
�"�l�Oف�J���C	��h��D���
�g�d�u�8�3���P���F�N����
� �g�`��l�K�������T��A�����0�<�0�&�0�8�_����ԓ�l ��X�*��y�c�|�_�w�}�W�������9��h\�B���u�h�&�1�;�:��������A��M�����1�%��9�����A����J��G����u�u�u�8��h����O�ѓ�F���*���<�
�0�!�%�/����Q����V��h8��G���d�
� �g�`��D��O����9F�N��U���
�c�3�
�a�l����Dӕ��l
��^�����'�'�&�/��4����	����9��h��G��
�f�y�c�~�W�W���Y����^��1��*��`�%�u�h�$�9��������G	��E�����<�;�1�<��8����M����O��=N��U���
�
� �d�o��F��Y����_	��T1�����}�0�<�0�"�.����Q����^��V�����e�g�%�|�b�t�L���YӒ��l_��Q��M���%�u�h�&�3�1��������AN��D��]���<�;�1�$��.����N����^��h�Y��|�_�u�u�:��F���&����l��S�����<�;�<�
��(�E��&����\��G1�����9�d�d�n�w�}����@����lT��1��U��}�8�
�a��8�(��HӞ����T�����d�d�n�u�w�)���&����
P��G\��H���<�;�<�
��8�(��IӞ����T�����d�d�n�u�w�)���&����S��G_��Hʦ�1�9�2�6�!�>����������^	��¤�
�&�<�;�n�;�(��A����U��UךU���8�
�`�3��m�G���Y���]��^	�����
� �f�c��n��������]��[��D��u�u�!�%�n����Iǹ��Z���*���
�0�
�d�c�%�Ͽ�&����G9��1�N���u�!�%�l��(�D��&���F��^	�����
�0�
�e�d�%�Ͽ�&����G9��1�N���u�!�%�l��(�D��&���F��h �����'�
�f�
�"�n�Eށ�K����W	��C��\�ߊu�u�8�
�n�;�(��I����[�L�����}��6�
�6�8�$�������lW��h��*��g�h�4�
�8�.�(���&����_��^�����u�8�
�
�"�l�Nށ�K���@��[�����6�:�}�=�1�����Q����V��V ��*���d�f�
�f�{�2��������]��Y��R��s�!�%�m�1��G���	����W��X����|�|�n�u�w�)����&����l��S�����:�&�
�#��}�W���&�Փ�V�� X�N���u�!�%�&�1��G���	�����h�����0�!�'�&�0�8�_�������l
��1��4���u�<�;�1������N���l�N��*����&�
�!�"�)����M˹��lT��1��U��_�u�u�u�w�8�(���LĹ��lT��1��U���;�}�'�6�9����HŹ��V�
N��R���9�0�_�u�w�}�W���&����9��h\�E���n�u�u� �#�;�(��N����[�L�����}�;�<�;�3�;����*����l'��X�����9�0�l�
��(�E��&���F��D�����-�
��-�"���������R
��hW��D���
�f�l�%�~�}����[����F�B �����"�d�3�
�o�m����D�ο�T��D�����3�
�m�g�'�}��������VW��h�����m�a�%�|�]�}�W�������D9��Q��G���%�u�h�}�:�n�N�������]9��h\�F���u�:�u�<�9�4�(���K����CU�=N��U���0�3�:�
��2�(���K����CT�
N����
� �g�m��o����&�ޓ�l ��\�*��n�u�u� �3�/����J����_��h�I���&�2�7�!�f�/���M�ƭ�WF��G_�����l�`�%�|�]�}�W�������D9��Y�����e�m�%�u�j�u���&����V��G\��ʥ�f�
�d�3��d�B���P���F��S�����a�3�
�d�g�-�W��Q����Q��1����l�u�;�u�:�l�(���J����CT�=N��U���0�3�:�
��2�(���J����CT�
N����
� �f�m��o����&�ޓ�9��h]�F���|�_�u�u�9�8����&����T��G\��H���<�;�4�&�0����A�����������d�d�<�3��m�D���P���WF��_��