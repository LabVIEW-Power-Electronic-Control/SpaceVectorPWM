-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǑ[�������n� �2��2�������T��_�[���n� �0���s�"���0����wH��[Uװ���!�u�c�����������G	��D��*���d�<�_�0�2�4�W�ԜY�ƅ�F�N��U���o�;�0�0�w�`�G�ԜY�Ƃ�~9��v)��U���o�;�0�0�w�`�F�ԜY�ƨ�]W��~*��U���u�u�<�!�0�/�M���K���F��Y\��<���u�u�u�u�>�)����C����l�N��ي���u�u�w�}�������F��d��Uʱ�;�
���w�}�W�������V�
N�N���u�1� �
��	�W���Y���Z��P��O���g�n�%�'�w�W�W������\��N�����2�6�#�6�8�u�FϺ�����O��N�����u�u�<�u�$�9��������G	��_�����:�e�n�u�w�9����Yɏ����h�����0�!�'�f�w�2����I��ƹF��^ �U���;�u�!�
�8�4�(��������Y��E��u�u�1� �w�}�Wձ�ӕ��l
��^�����'�f�u�:�9�2�G���s����V��C����=�!�6� �2�/�ϱ�Y����v$��r��*���
�!�d�&�;��E�����F���ʼ�!�'�4�u�>�3��ԜY�ƿ�T����U���o�&�1�9�0�>��������W	��C��\�ߊu�u�x�9�!�1�Fϭ�����9F������8�-�d�e�w�}�W���&����P9��T��]��1�"�!�u�~�W�W���������h_��U���o�&�1�9�0�>����������Y��E��u�u�x�u�2�8�W�������@l�N�����u� �
�
�w�}�Mϭ�����Z��R����u�:�;�:�g�f�������_F�
��A�ߠx�u�0�0�6�8��������\��=��*ۊ�u�h�1�;�w�5�ϭ����F�N�����<�g�_� ���W������9l�)�����0�9�#�9�e�1��������lV�
N�����e�"�0�u�2�u�^��^����_��Z��D��_�x�u� �'�)��������GF���*؊�n�_�;�u�%�5��������