-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ������}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e���o��}�#���6����e#��x<��F���:�;�:�e�l�}�WϿ�&���/��d:��9����_�u�u���(���	����\��yN��1�����_�u�w��(���&����z(��c*��:���
�����l��������l�N��D���-��4�
�;�}�W���*����|!��d��Uʥ�g��'�:�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����c��X
�����1�o��u���8���B�����h;�����2�0�e�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���&ǹ��g��Y	��*ڊ�%�#�1�o��	�$���5����l�N��A����8�;�
��}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y����lR��h:�����0�d�4�
�;�}�W���Y����)��tUךU���
�
�
�u�w��$���5����l0��c!��]��1�"�!�u�~�W�W���&ƹ��e9��h��U���������}���Y����e9��Z��*���u�u� �u���8���&����|4�_�����:�e�n�u�w�-�A���-����T9��1��*���u�u� �u���8���B�����h8�����2�0�d�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���&Ź��g��Y	��*ۊ�%�#�1�o��	�$���5����l�N��B����o��u���8���&����|4�_�����:�e�n�u�w�-�@���/����E
��N��U���
���n�w�}����.����Z��R1�Oʚ�������!���6���F��@ ��U���_�u�u�
����������l��A��Oʚ�������}���Y����d9��Z��*���u�u� �u���8���&����|4�_�����:�e�n�u�w�-�O�������T9��1��*���u�u� �u���8���B�����1�����u�u� �u���8���&����|4� N�����u�|�_�u�w��B�������R��[
��U���u��
���}�L����ƓR��^�����u�0�4�u�1�0�5���<����F��d��Uʴ�!�<� �0���(���<����|(��y(��Oʆ���n�u�w�<��������|4��p+��'����
���8�}����Y�ƭ�P��R�����&�u�u�w�b��4�������_��G1�Dފ�y�����	�#���D����{*��~ ��!�����e����'���?����W��{=��;���
���-�`�m�G���M���.��h'�� �����h�`�g�m�G���5����c3��v<��H���0�&�����4���2����V��^��9����
��h�c��$���7������RB��&������e���$���=���.��h=��*���d�a�y����(���D����ND��N�����!�;�u�%�4�3��������\��c*��:���u�h�r�r�]�}�W���
������T�����2�6�e�o���;���:���V�=N��U���&�4�!�4��	��������\��c*��:���
�����}�������	[�^�E���_�u�u�:�$�<�Ͽ�&����GT��D��U����
�����#���Q�ƨ�D��^��O���e�e�d�w�]�}�W���
������d:��ي�&�
�u�u���8���&����|4�N�����u�|�o�u�g�m�G���s���P	��C��U����
�!�
�$��W���-����t/��a+��:���`�1�"�!�w�t�M���I����D��N�����!�;�u�%���ځ�
����	F��s1��2������u�b�9� ���Y���F�^�E��u�u�6�;�#�3�W���*����9��Z1�Oʆ�������8���Lӂ��]��G��H���e�e�e�n�w�}��������R��X ��*���g�e�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�e�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�f�f�W�������R��V�����
�#�g�d�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�g�l�L���YӅ��@��CN��*���&�
�#�g�e�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����\��V �����:�&�
�#�e�n�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��B�����D��ʴ�
�:�&�
�!�o�C��*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��X �����4�
�:�&��+�(���Y����)��t1��6���u�e�1�"�#�}�^��Y���9F������!�4�
�:�$�����L����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����4�!�4�
�8�.�(���&����`2��{!��6�����u�d�3�*����P���V��d��Uʶ�;�!�;�u�'�>��������
U��[��Oʆ�������8���O�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��d�e�e�d�f�m�F��I����V��_�N���u�6�;�!�9�}��������EP��[�@���u�u��
���(���-���U��X����u�h�w�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�D��d�e�n�u�w�>�����ƭ�l��D�����f�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��d�d�d�w�]�}�W���
������T�����f�
��o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�d�d�g�f�W�������R��V�����
�#�g�d�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�f�m�U�ԜY�Ư�]��Y�����;�!�9�f���Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�l�G��B�����D��ʴ�
�:�&�
�!�o�F���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��H����F�T�����u�%�6�;�#�1�E؁�Y�Ɵ�w9��p'��#����u�g�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��B�����D��ʴ�
�:�&�
�!�o�F���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��H����F�T�����u�%�6�;�#�1�D݁�?����u �=��*����
����u�FϺ�����O�
N��D��d�d�d�d�f�l�F��H����W��_�����u�:�&�4�#�<�(���
���� T��^�E��o������!���6���F��@ ��U���o�u�d�e�g�m�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D�����g�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��d�e�e�w�]�}�W���
������T�����f�
�u�u���8���&����|4�^�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�f��}���Y����G�������!�9�g�d�m��3���>����v%��eN��U���;�:�e�u�j��F��Y����\��V �����:�&�
�#��}�W���&����p9��t:��U��1�"�!�u�~�g�W��H����F�T�����u�%�6�;�#�1�C��Cӵ��l*��~-��0����}�u�:�9�2�G���D����V�=N��U���&�4�!�4��2�����ԓ�u ��q(��Oʆ�������8���J�ƨ�D��^��O���d�d�d�d�f�l�F��H����W��_�D��n�_�u�u�>�3�Ͽ�&����@�=��*����
����u�W������F��L�E��w�_�u�u�#�/����Y����V��S��U���!�<�2�_�w�}��������U��R �����u�3�4�
��;���
����_F��L�����_�u�u�<�9�1��������V��c1��D���8�e�o����0���s���@��V�����2�7�1�g�w�}�8���8��ƹF��^	��ʥ�e���<��4�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1��4���%�0�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�u�W�W���������h/��*���#�1�<�
�>�}�W���&����p]ǻN�����9�%�e���<�(���&����\��c*��:���u�h�r�r�]�}�W�������lW��V��*���&�2�o����0���/����aF�N�����u�|�_�u�w�4����	�ד�R��h����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�n�u�u�$�:����&¹��K9��V�����;�&�2�o���;���:���F��P ��U���
�4�
�
�'�+��������`2��{!��6��u�e�n�u�w�.����Y����c��X
�����2�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�K����Z	��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�>�3�Ϯ�K����Z	��V�����;�&�2�o���;���:���F��P ��U���
�0�<�1�6��������5��h"��<���h�r�r�_�w�}����Ӗ��l$��h�����o������!���6���F��@ ��U���_�u�u�<�9�1����;����A��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�&�2�4�w��(���&����_��Y1���������W�W���������h,��*���#�1�%�0�w�}�#���6����	[�I�U���&�2�4�u���(�������\��c*��:���
�����l��������l�N�����u�
�
�
��/���*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��^	��ʥ�b���4��1�(���
���5��h"��<��u�u�&�2�6�}�(؁�&����l��h���������g�W��B�����Y�����<�
�1�
�g�}�W���5����9F������&�2�7�!�%�:�N��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��#���
�
�0�
�g�i�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��Z��B���2�d�e�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӗ��R��P ��*���f�b�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӗ��R��P ��*���
�e�`�o���;���:����g)��^�����:�e�n�u�w�.����Y����9��hZ�*��o������!���6��� F��@ ��U���_�u�u�<�9�1����M����lW��N�&���������W��Y����G	�UךU���<�;�9�3�'�3�������� 9��Q��AҊ�f�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�	����V9��E��F���'�2�d�g�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����R��^	������
�!�
�$��W���-����t/��=N��U���;�9�4�
�>�����J����q)��r/�����u�<�;�9�'��݁�L����W��G\��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u��<�E��&����V��T��!�����
����_������\F��d��Uʦ�2�4�u�8��n����H����	F��s1��2������u�g�9� ���Y����F�D�����8�
�g�<�1��Eف�K����g"��x)��*�����}�u�8�3���B�����Y�����d�
�
�0��m�G��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��G1��؊�
� �c�c�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��a��*���0�
�e�`�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������C9��P1������&�f�3�:�o�Mύ�=����z%��N�����4�u�%�&�0�?���O����|)��v �U���&�2�4�u�/���������`0��U��%���6�<�&�'�0�l�B���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*���
�&�$���)�(���&����`2��{!��6�ߊu�u�<�;�;�<�(���&����S��N��:����_�u�u�>�3�Ϲ�	����l ��h��G���4�
�:�0�m��3���>����F�D�����-�
�:�0�#�/�(�������c9��T��D���2�d�`�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�C9��S�������7���.����K����lW��N�&���������W��Y����G	�UךU���<�;�9� ��2��������~��q6�����<�d�'�2�f�k�W���-����t/��a+��:���b�1�"�!�w�t�}���Y����R
��g_��*���c�e�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƃ�9��E��D��u�u��
���(���-���U��X����n�u�u�&�0�<�W�������A9��X��D���
�c�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƥ�l
��q��9���
�d�'�2�f�j�W���-����t/��a+��:���d�1�"�!�w�t�}���Y����R
��G1�����0�
��&�b�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������U�� [��G��������4���Y����\��XN�N���u�&�2�4�w�8�(���&����T9��]��U���
���
��	�%���Y����G	�UךU���<�;�9�0�>�>����&����U��N�&���������W������\F��d��Uʦ�2�4�u�0��0�E�������9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�(�������
W�=��*����
����u�W������]ǻN�����9�2�%�3��m�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����!�g�'�2�f�m�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h8��G���
�0�
�d�o�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������C1�����d�d�u�u���8���&����|4�N�����u�|�_�u�w�4��������9��P1�D���u��
����2���+����W	��C��\�ߊu�u�<�;�;�/����˹��lQ��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u���(�������T��N��1��������}�GϺ�����O��N�����4�u�4�2�f�<��������U��[��G��������4���Y����\��XN�N���u�&�2�4�w�<��������]��1����g�u�u����>���<����N��S�����|�_�u�u�>�3�ό�����R
��M�����
�b�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���:�
�0�
�f�i�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��E1��*���
�:�%�d���(߁�&����W��N�&���������W��Y����G	�UךU���<�;�9�4��4�(�������@��Q��@�������W�W���������D�����g�e�o����9�ԜY�ƿ�T����*����'��:��d�E���I�Փ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���?����\	��W��*���
�
� �l�e�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�f��(���&¹��l_��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�6�/��������\��1�����f�3�
�c��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�����'��:�
�n�o����L����
Q��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%��(߁�&����lT��h�����!�o�����4�ԜY�ƿ�T��	��*���
�
�
� �e�n�������5��h"��<��u�u�&�2�6�}����&ù�� 9��h\�*���'�4�,�o���;���:���F��P ��U���
�
�
�
��(�E�������C��1��Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-�����Փ�F9��1��*���
�
�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U9��Q1�����l�
�;�7�#��(���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����e�3�f�3��d�(�������]9��N��1��������}�D�������V�=N��U���;�9�2�%�1�m�������� 9��h�� ���d�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����l ��h��G���4�
�0� �9�o�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E��*ڊ�
�
� �g�d�<�(�������\��c*��:���
�����}�������9F������2�%�3�e�1�n����@����l��N��1�����_�u�w�4��������w#��e<�����c�0�e�'�0�o�D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����<�����!�'��i��������P�=��*����
����u�FϺ�����O��N�����4�u�'�
�#���������lT��h^��*���
�g�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����_��X�����d�
�
�
��8�(��Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y���������2�0�Cہ�&¹��T9��N�&���������W��Y����G	�UךU���<�;�9�6���2���+����lR��R1�����g�m�o����0���/����aF�N�����u�|�_�u�w�4��������l ��h"�����'�2�g�d�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƫ�C9��1��F���
�l�
�%�$�<����&����G9��PN�&������o�w�m�L���Yӕ��]��P�����e�
�e�o���;���:����g)��]����!�u�|�_�w�}����ө��l0��h�����
�f�
�d�m��3���>����v%��eN��Eʱ�"�!�u�|�]�}�W�������cW��h_��*���`�c�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƃ�9��Q��Eڊ�d�o�����4���:����P��S�����|�_�u�u�>�3�Ϲ�	���� V��G_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%����I����	F��s1��2������u�a�}�������9F������!�%�<�3��l�(��Cӵ��l*��~-��0����}�g�1� �)�W���s���@��V�����
�
� �f�o�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��E1�����g�
�g�o���;���:����g)��]����!�u�|�_�w�}����ӕ��]��h��F���%�u�u����>���<����N��
�����e�n�u�u�$�:����&����lP��B1�B���u�u��
���(���-���V��X����n�u�u�&�0�<�W������� S��G_��U���
���
��	�%���Iӂ��]��G�U���&�2�4�u�:��A���&����CV�=��*����
����u�GϺ�����O��N�����4�u�8�
�a�;�(��&���5��h"��<������}�a�9� ���Y����F�D�����8�
�b�3��j�(��Cӵ��l*��~-��0����}�e�1� �)�W���s���@��V�����m�3�
�m��l�Mύ�=����z%��r-��'���e�1�"�!�w�t�}���Y����R
��Z��M���
�m�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƾ�U��W��G��������4���Y����\��XN�N���u�&�2�4�w��(���&����
W��N�&���������W������\F��d��Uʦ�2�4�u�7�#�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʥ��9�
�d�1��Eׁ�K����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
� �c�n����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��#���3�
�e�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������hY��*���a�f�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��^1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������l��B1�B���u�u��
���(���-��� W��X����n�u�u�&�0�<�W����ԓ�l ��]�����u��
����2���+������Y��E��u�u�&�2�6�}��������l ��]�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)��������R��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�%��.����&����G9��hZ�*��o������!���6�����Y��E��u�u�&�2�6�}��������Z9��hZ�*��o������!���6�����Y��E��u�u�&�2�6�}����&����_��N�&���������W������\F��d��Uʦ�2�4�u�0�2�8�(�������lR��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��2�(���&����V��N�&���������W������\F��d��Uʦ�2�4�u�'�2�:�(���&����P��N�&���������W������\F��d��Uʦ�2�4�u�8���D���&����CT�=��*����
����u�W������]ǻN�����9�%�f�
�����L����	F��s1��2������u�g�9� ���Y����F�D�����'�0�2�a��8��������l ��W�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)��������]9��h[�*��o������!���6�����Y��E��u�u�&�2�6�}��������U��W��G��������4���Y����\��XN�N���u�&�2�4�w�+��������_��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�m����Kù��\��c*��:���
�����}�������9F������7�8�'�0�>�4����&����CT�=��*����
����u�W������]ǻN�����9� �1�'�;�*��������T��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�%��1�(ځ�����U��\��F��������4���Y����W	��C��\�ߊu�u�<�;�;�-�!���&ƹ��U��^��F��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����^��N�&���������W��Y����G	�UךU���<�;�9�!�'�j�(���L�ޓ� F��d:��9�������w�m��������l�N�����u�
�
� �b�o����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���<�3�
�l��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��^��*���`�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӗ��R��P ��*���c�g�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӗ��R
��Z�� ���e�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����W��h��C���%�u�u����>���<����N��
�����e�n�u�u�$�:��������\��h��C���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϱ�&����R��D�����
�m�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������K��C1�����:�
�c��1��N܁�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�c�3�
�e��F��*����|!��h8��!���}�c�1�"�#�}�^�ԜY�ƿ�T����*���3�
�a�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����A9��Q��G݊�g�o�����4���:����V��X����n�u�u�&�0�<�W�������lT��^1��*���
�a�o����0���/����aF�
�����e�n�u�u�$�:��������Z��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������l��B1�D���u�u��
���(���-��� W��X����n�u�u�&�0�<�W����ԓ�
9��hY�*��o������!���6���F��@ ��U���_�u�u�<�9�1����Nʹ��lQ��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��G�������9��T��!�����
����_�������V�=N��U���;�9�6�'�.�o����Iǹ��\��c*��:���
�����}�������9F������%�f�
�
�f�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�c�
�
�"�e�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����0�
�0�:�����@����	F��s1��2������u�g�9� ���Y����F�D�����<�;�<�
�8��(���A�Г�F��d:��9�������w�m��������l�N�����u�
�l�1�:�/����&����l^��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2���������U��_��G��������4���Y����\��XN�N���u�&�2�4�w��N�������]9��Y�����
�`�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ʈ�^��R1�����!�<�3�
�c��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��Y�����3�
�g�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����Q��E	�����
�`�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƽ�e��h\�*���
�
� �m�b�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1��؊�
� �m�f�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��a��*���3�
�m�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������O=�����
� �!�4�#�n�(���A�ߓ�F��d:��9�������w�n�W������]ǻN�����9�4�'�9��2�(���	����9��1��*��
�a�o����0���/����aF�N�����u�|�_�u�w�4��������G9��E1�����l�e�0�e�e�;�(��&���5��h"��<������}�f�9� ���Y����F�D�����'�
�!��%�����@�ԓ�lV��B1�A���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����\��X��Dӊ�
�
�
�
�"�d�O���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����9�
�:�
�8�-�Fց�&����U��V��G��������4���Y����W	��C��\�ߊu�u�<�;�;�<����&����	��h_��G���d�g�3�
�b��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*����'��:��d�E���H�ғ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�-�9���
����`2��{!��6�����u�`�3�*����P���F��P ��U���&�2�7�1�f�o�MϜ�6����l�N�����u�%�&�2�5�9�C���Y����v'��=N��U���;�9�4�
�>�����J����q)��r/�����u�<�;�9�6���������\��x!��4��u�u�&�2�6�}��������lS��N��:����_�u�u�>�3�Ͽ�&����Q�� _��U�����n�u�w�.����Y����Z��S
��A������]�}�WϽ�����]��,��6���3�e�3�f��W�W������9F�N��U���6�>�o��w�	�(���0��ƹF�N�����!�o��u���8���B���F������!�o��u���8���B���F������u�u� �u���8���B���F������u�u� �u���8���B���F������,�o�����;���:���F�N��*���=�
�
�u�w��$���5����l0��c!��]��1�"�!�u�~�W�W���Y�ƥ�l��h\��U���������!���6���F��@ ��U���_�u�u�u�w�3����&ù��	F��=��*����
����u�FϺ�����O��N��U���4�
�0� �9�m�Mϑ�-ӵ��l*��~-��0����}�d�1� �)�W���s���F�V�����;�d�o����3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���Y����V��Y1�Oʚ�������!���6���F��@ ��U���_�u�u�u�w�-��������	F��cN��1��������}�@Ϻ�����O��N��U���4�
�0�o��}�#���6����]ǻN�����:�%�;�;�l�W�}������F��G1��E���f�3�
�l�w�}��������^S��q-��6���
�
�_�u�w�2�ϳ�	��ƹF�N�����>�h�u�%�4�6�}���Y���R��D��Kʴ�
�&�y�u�w�}�WϿ�&����GF�	��*���
�
�
� �e�n��������9F�N��U���1�;�u�k�0�-�����Փ�F9��1��*���0�_�u�u�w�}���������h��*���
� �g�f�6�����s���F�V�����u�k�2�%�1�m�������� 9��h�����u�u�u�u�>�����&¹��X��E��*ڊ�
�
� �g�d�4�(�������eJǻN��U���;�8�-�g��`�W���&����U9��Q��Lي�;�8�-�g��W�W���Y�ƥ�l��V1��#��u�'�
�
���(���K�Փ�]9��C��*���u�u�u�u�6��������F��G1��E���f�3�
�l��-��������9F�N��U���'�!�'�
�w�c�����֓�lU��B1�F���
�0� �;�f�W�W���Y�ƭ�l��B��G��u�'�
�
���(���K�Փ�C9��C��*���u�u�u�u�6��������F��G1��E���f�3�
�l��-��������9F�N��U���6�u�k�2�'�;�G���J����_��V����_�_�_�u�w�p��������]��C��U´�
��3�8�w�;����
������_��[���_�u�u�%������
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��h-�����i�u�%���)�(���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�V�N��U���u�u�u�u�w�}����*����Z�V��&���8�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��E��*ڊ�
�
� �g�d�<�(�������l��E�����&�<�;�%�8�8����T�����h��*���
� �g�f�6�����&����G��h��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�'���(���&����
U��G1�����4�
�!�'��8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�d�;���P�Ƹ�V�N��U���u�u�u�u�w�}�����֓�lU��B1�F���
�!�'�
�'�.�������F��h�����:�<�
�n�w�}�W���Y���F��[��U���%�6�;�!�;�:���DӁ��l ��h��*���g�f�4�
�2�9�^������F�N��U���u�u�u�u�0�-�����Փ�F9��1��*���'�
�%�&�6�)����E�ƭ�l��D�����
�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��4���4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�e���<�(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�
�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����4�
�<�
�3��D�������9F�N��U���u�u�u�u�w�}�W���&����R��[
�����i�u�%�6�9�)��������F�N��U���u�u�u�u�2�.����	����l��hZ�U���;�_�u�u�w�}�W���Y���F�N��E����4�
�9��/���Y����r9��V����u�u�u�u�w�}�W���Y����]��QUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�֓�l0��E�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��a1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���(������F��h�����#�g�e�_�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���
�
�
�%�!�9�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�|�u�?�3�}���Y���F�N��U���%�e���'�8�W��	�֓�l0��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����e9��h��*���2�4�&�2�w�/����W���F�G1������4�
�9��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h��*���%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��F��*���
�1�
�f�~�)����Y���F�N��U���u�u�u�u������&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lR�����ߊu�u�u�u�w�}�W���Y���F��1�����4�
�9�
�%�:�K���&¹��K9��V����u�u�u�u�w�}�W���Y����]��QUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ד�R��h��ʴ�&�2�u�'�4�.�Y��s���C9��Z��#���0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(ށ�����C��R�����:�&�
�#�e�m�}���Y���F�R�����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t���������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*ۊ�4�
�
�%�!�9�^������F�N��U���u�u�u�u�'�l����/����TF���*���
�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��%���:�
�%�#�3�-����
������T��[���_�u�u�
��8��������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�2�4����&����C��R�����:�&�
�:�>��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�3��-�������� _�C��U���u�u�u�u�w�}�W���Y�����h>�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�m�w�5��ԜY���F�N��U���u�u�u�%�e�����&����_��E��I���
�
�0�<�3�<�(���B���F�N��U���u�u�u�;�w�;�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u�
�
�0�>�9����Y����T��E�����x�_�u�u����������T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�g��'�:��/���Y����\��h��G��_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ԓ�V��S1��*���|�|�!�0�w�}�W���Y���F�N��U���
�0�<�1�'�8�W��	�ԓ�V��SUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ӓ�l0��G1�����0�u�&�<�9�-����
���9F���*���
�%�#�1�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��u1�����9�
�'�2�k�}��������\��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����UF��G1�����1�b�l�u�?�3�}���Y���F�N��U���u�u�%�`����������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&���G��d��U���u�u�u�u�w�}�W���YӖ��l$��h�����%�0�u�h�'�h�5�������W]ǻN��U���u�u�u�u�w�}�������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u���(�������@��YN�����&�u�x�u�w�-�B���/����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�`���%�2�}�JϿ�&����G9��\��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��h[��*���'�2�i�u���(��Y���F�N��U���;�u�3�u�w�}�W���Y����]��QUךU���u�u�;�u�1�W�W����Ƽ�\��DUװ���u�x�%�b����������V��D��ʥ�:�0�&�u�z�}�WϮ�N����l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}��������W9��G�����_�u�u�u�w�}�W���Y���F�G1��6���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�a�w�5��ԜY���F�N��U���u�u�u�%�`��!���&����C��R�������4�
�;�f�W���Y���F�N��U���;�u�3�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*݊�
�
�'�2�6�.��������@H�d��Uʥ�b���%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��a1�����h�4�
�:�$�����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�<����	����@��X	��*���u�
�
�
��-����P�Ƹ�V�N��U���u�u�u�u�w�}����:����A��S��*݊�
�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�^"�����'��:�
��8�(��Y����T��E�����x�_�u�u��1�(���&����l��R	��Mۊ�&�<�;�%�8�}�W���������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�P���Y����9F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��C���8�`�|�!�2�}�W���Y���F�N��U����9�
�:��2��������W�
N��*����'��:��l����H����9F�N��U���u�u�u�9�>�}��������W9��G�����_�u�u�u�w�}�W���Y���Z*��^1�����:�
�
�0��e�W������]��[��E�ߊu�u�u�u�w�}�W����ƥ�l�N��U���u�0�1�<�l�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�W���T�ƭ�@�������{�x�_�u�w�/����Yۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�p�z�W������F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�a�3�:�n�W���Y������T�����2�6�e�h�0�-�����Փ�F9��1��*���0�|�|�!�2�W�W���Y���F�N��D���'�2�d�b��t�K���)¹��U��^��D��n�u�u��f�����H����O�
N��D���3�
�c�
�f�l�L���Yө��l0��R	��E��g�u�h��f�����Où��T�=N��U���
�
�0�
�g�m�D���Dө��l0��B1�E���}�|�_�u�w��(�������V�N�U���
�
� �c�g�-�_���s���|6��a1����b�}�|�i�w��(�������l��G�U����d��'�0�l�@���P���|6��a1��*��
�d�c�n�w�}�8���/����lW��F�U���d��3��k�(��N��ƹF��g_��*���
�e�e�m�w�`�8���/����P��G_��\�ߊu�u��
��8�(��I���[��g_��*���c�e�%�}�~�W�W���)¹��A��^�]��u�h��d��;�(��&���O��N��:����'�2�d�`�u�F���Dө��l0��B1�E���}�d�n�u�w��F�������Q��\��I����
�
� �a�m����K��ƹF��g_��*���
�e�e�d�~�a�W���&����lP��h�D���_�u�u�������I���O�
N��D���3�
�c�
�f�l�^�ԜY�ƃ�9��E��D��}�`�u�h��l�!���&����CW�G�U����d��'�0�l�@���O���)��h8�� ��e�%�}�c�l�}�Wϑ�H����V��Y�D���i�u��
��(�A���	����]ǻN��%ۊ�
�0�
�e�g�l�^��Y����e9��hX�*��d�|�_�u�w��(�������V�G��Hʚ�d��3�
�a��F��P���F��1�����d�b�}�e�w�`�8���/����P��G_��E��u�u��d��/���N����F�!��*��� �c�e�%��l�L���Yө��l0��R	��E��g�|�i�u���(���O�֓�N��UךU����
�
�0��m�G��P���|6��a1��*��
�d�g�|�]�}�W���&����T9�� ^��A���h��d��1��A߁�H����l�N��D���'�2�d�b��h�W��6�ד�l ��X�����`�n�u�u��l�!�������N��N�U���
�
� �c�g�-�_��B���)��h8�����e�e�g�|�k�}�'ށ�&����V��F�\�ߊu�u��
��8�(��I����Z�x>��#���
�c�
�d�e�t�}���Y����e9��P1�B���l�u�h��f�����Où��T��d��Uʚ�d��'�2�f�j�_��Y����cW��h��C���%�}�e�n�w�}�8���/����lW��F�\��u��
�
�"�k�G���Q���9F�N��U���u�u�u�-��2��������~��q6�����<�d�'�2�f�h�W������lV��h]�� ��f�4�
�0�"�3�F�ԜY���F�N��Uʳ�%�;�1�
�2�0�$�������l��A��*���
�e�e�i�w�/�(���&����U��]�����!�'�
�n�w�}�W���Y���F��O�����!�'�
��6�>�/�������@9��P1�@���h�2�%�3�g�;�D���&����R��R����_�u�u�u�w�}�W���Y����\��C��*���4�6��
�%�+�(ށ�����S�
N�����e�3�f�3��d�(�������]9��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}���Y���R��P �����&�{�x�_�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�`�1�0�C�������K��X �����
�c�
�g�j�<�(���
����9��G�����u�u�u�u�w�}�W���+����9��[1�����
�0�
�d�o�a�W����ד�_
��Y��G���
�c�
�g�]�}�W���Y���F�e��ۊ�9�
�0�:��8�(��M���a��R_�����0�:�
� �`�l���Y���F�N��U���
�4�g�`��8�(��A���T��Q��Eڊ�g�`�u�:�9�2�E���s���F�N��U���$�<�
�
�2��F��E�ƫ�C9��h]�*��g�u�:�;�8�o�^�ԜY���F�N��Uʧ�<�<�<�
�2��F��E�ƾ�Z9��^V�� ��l�%�n�u�w�}�W���Y�����h��G���'�2�d�l�w�`��������Z9��hX�*��_�u�u�u�w�}�W���Y����G��^1����m�u�h�&�;�)��������9��d��U���u�u�u�u�w�.�����ԓ�V��^�I���'�
� �f�g�-�_������\F��UךU���u�u�u�u�w�}����N����lW��N�U���
� �f�e�'�u�NϺ�����_�=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}���Y���R��P �����&�{�x�_�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�c�1�0�B���Y����9F�N��U���u�u�u�'��)�1���5����_��h��*܊�0�
�g�u�j�<����&����	��h_��G���e�`�3�
�c��D�ԜY���F�N��Uʴ�'�9�
�:��2���&����9��P1�G��u�'�
�!��/�;���&�ߓ�l��h_�� ��l�%�n�u�w�}�W���Y�����~ ��-���!�'�
�a�2�m����K���F��E1��*���
�:�%�d���(߁�&���� S��UךU���u�u�u�u�w�}����=����a��Z1�*���
�0�
�`�w�`��������A9��X��L���0�d�f�3��k�(��s���F�N��U���6�
��������MŹ��9��P1�F��u�'�
�!��/�;���&�ߓ�l��h_�� ��d�%�n�u�w�}�W���Y�����~ ��-���!�'�
�c�2�l����K���F��E1��*���
�:�%�d���(ށ�&����Q��UךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��ԶY���F��D��U���6�&�{�x�]�}�W���������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�P���Y����9F�N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�e�;���P�Ƹ�VǻN��U���u�u�u�u�/���������U��h��*��`�i�u�-��2��������l0��B1�M���n�u�u�u�w�}�W���YӖ��R
��[�����e�e�i�u��<�E��&����T��UךU���u�u�u�u�w�}����K����V��Z�I���8�
�g�<�1��Eف�K���F�N��U���u�!�%�b��8�(��L���C9��[\��@���
�d�
�g�d�}��������l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�^Ϫ����F�N��U���u�<�
�<��/�;���&�ד�V��Y�I����9�
�:��2���&����_��UךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��ԶY���F��D��U���6�&�{�x�]�}�W���������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�P���Y����9F�N��U���u�3�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�d�j�<�(���Y����]	��V�����1�
�e�|�~�)��ԜY���F�N��Uʥ��9�
�
�2��G��E�Ƽ�e��hX�� ��b�%�}�l�3�*����A��ƹF�N��U���u�u�7�4�$�:�(ہ�����S�
N��*���<�;�a�3��d�(��s���F�N��U���'��a�'�0�l�E���DӔ��lR��B1�D���n�u�u�u�w�}�W���Yӕ��]��h��*��u�h�&�2�5�)����Jʹ��P��S�����e�n�u�u�w�}�W���Y����^�� 1����e�u�h�!�'�k�(���J�ӓ�N��
�����`�|�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=N��U���4�&�2�u�%�>���T���F��X�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������A��N���ߊu�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�Փ�@��G�����_�u�u�u�w�}�W���Y����_T��h��*��`�i�u�
�6�o����&����CU��N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�W���6�ד�l��h_�E��u�:�;�:�d�t�K���I����V��^�E��e�e�e�e�g�m�G��B���F���U���!�&�4�0��-�9���
����UF��RN�����8�6�<�0�w�p�W�������l ��h�����%�:�u�u�%�>��������l ��N��*���u�%�&�2�5�9�F��Y����U9��Q1�����l�
�%�1�9�q��������Z9��hX�*��_�u�u�0�>�W�W���Y�Ư�@��G1��*���u�&�u�u�w�}�W�������R��c1��D���8�e�h�u�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN��´�
�<�
�1��m�^�������F�N��U���u�u�u�u�6��$������R��c1��G���8�d�_�u�w�}�W���Y���V
��=N��U���u�u�u�u�w�}�W���7����^F���&���!�
�&�
�l�}�W���Y���F���U���_�u�u�u�w�}�W���Ӈ��`2��C\�����u�k�_�u�w�}�W���Y���R��d1����u�%��
�#�����B���F�N��U���;�4�
��$�n����K���9F�N��U���u�u�u�%������DӇ��`2��CZ�����n�u�u�u�w�}�Wϩ��ƭ�l5��D�����f�h�u�u�w�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R��Y��]���6�;�!�9�0�>�G������lV��h]�� ��f�4�
�:�2�t�^Ϫ����F�N��U���u�u�u�4������E�ƭ�l5��D�����a�_�u�u�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}��������l��h��*���k�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ����F�����;�
�
� �a�n����Y����\��h��*���|�u�=�;�w�}�W���Y���F�N�����
�&�u�h�6��#���H����lV��N��U���u�u�u�u�2�.�}���Y���F�N��U���4�
��3�:�a�W���*����9��Z1����u�u�u�u�w�}�W���Y����F�N��U���"�0�u�%���ف�
����X�N��U���u�u�u�u�6��$������R��c1��@���8�a�_�u�w�}�W���Y����	��R��H���_�u�u�u�w�}�W���Y����`9��ZN�Uȍ���w�_�w�}�W����Ư�@��N�����%�:�0�&�]�}�W���Y����e9��^1��*���
�d�i�u�#�����&����\��R��¦�2�0�}�
������I���R�dךU����
�
� �a�m����Dӕ��l
��^�����'�'�&�/��3����ۖ��l6��^�����<�|�c�|�l�}�W���Yө��l0��B1�E���u�h�&�1�;�:��������A��M�����1�3�%�9��2�(���	����e9��hX�*��y�a�|�_�w�}�W���6�ԓ�l��V�����f�
�d�i�w�)�(�������P�������&�2�0�}�����K����P��UװU����;�0�
�;�����K����P��G\��H���w�"�0�u�'�����&�ѓ�l �� [�����u�%�6�;�#�1�C���Y����D��d��Uʇ�;�0�
�9��8��������l��S��D���=�;�}�
�2�(���&����lQ��h�Hʴ�
�:�&�
�!��^ϻ�
���]ǑN��X���%�1�;�u�$�4�Ϯ�����F�=N��U���1�;�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
�ӓ�@��N�����;�
�
� �a�n����Y����V��=N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�b�;���Y����]	�������1�<�3�
�a��E������]��[��E���|�!�0�u�w�}�W���Y����C9��Y��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����VF��D��U���6�&�{�x�]�}�W�������R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�}���Y����]l�N��Uʼ�u�}�:�}�6�����&����P9��
N��*���'�|�u�;�w�<�(���
����T��N�����<�
�&�$���ށ�
����O��_�����u�u�u�u�w�-����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�1�0�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�4�
�2�9�W�������A	��D�X�ߊu�u�%�'�6�$��������\������}�%�6�y�6�����
����g9��1����u�-�!�:�3�4����O����l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����0�<�6�;�����J����F��h�����#�
�|�|�w�5��ԜY���F�N��*���1�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����V��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����1�d�c�4�$�:�W�������K��N�����<�
�1�
�g���������PF��G�����4�
�!�'�{�-�G���/����E
��^ �����%�d�8�-��<�(���&����Z�G1��%���:�
�%�#�3�4�(���UӖ��l$��h�����<�
�<�y�'�j�4�������W9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�d�c�i�w�u�(؁�&����l��h�����h�4�
�:�$�����&����AF��h[��*���%�#�1�<��4�W���	����@��X	��*���:�u�%�g��/����	����l��D��Hʴ�
�:�&�
�8�4�(�������lW��V��*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�e���<�(���&����Z������!�9�2�6�g�}����	����A������!�9�2�6�g�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����u�:�;�:�f�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����u�:�;�:�e�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*���u�h�}�%�4�3����H�����t=�����u�:�;�:�d�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����l��F1��*���
�&�
�y�0�-�����Փ�F9��1��*���0�_�u�u�2�4�}���Y���F�N�����<�
�1�
�a�}�J�������]��[����h�4�
�<��.����&����U��G�����:�}�4�
�8�.�(�������F��G1��E���f�3�
�l��-����P����F�R �����0�&�_�_�w�}�ZϿ�&����Q��Y����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h-�����_�u�u�0�>�W�W���Y���F�N��*���
�1�
�b�w�`�_�������l
��h_��U����
�&�}�w�2����M����F�R �����0�&�_�_�w�}�ZϿ�&����Q��_����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h-�����_�u�u�0�>�W�W���Y���F�N��*���
�1�
�d�w�`�_�������l
��h_��U����
�&�}�w�2����L����F�R �����0�&�_�_�w�}�ZϿ�&����Q��\�����;�%�:�0�$�}�Z���YӇ��@��U
��G؊�&�<�;�%�8�}�W�������R��d1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�g�i�w�<�(��������Y��E���u�%�6�;�#�1�F��B����������n�_�u�u�z�}��������lR��V�����'�6�&�{�z�W�W���	����l��hZ�����2�
�'�6�m�-����
ۇ��@��CB�����2�6�0�
��.�F������C9��v1�����9�|�u�u�5�:����Y���F�N��U���&�2�7�1�c�}�J�������]��[����h�%�e���<�(���PӇ����F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�u�9�}��������_	��T1�Hʴ�
�!�'�|�~�f�W�������A	��D����u�x�u�%�$�:����M�ƭ�@�������{�x�_�u�w�-��������
9��D��*���6�o�%�:�2�.����������D�����
��&�d�1�0�G���&¹��K9��V�����u�u�7�2�9�}�W���Y���F������7�1�a�u�j�u����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����4�
�9�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���Y����T��E�����x�_�u�u�'�.��������R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����\��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�m�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h>�����4�
�9�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���Y����T��E�����x�_�u�u�'�.��������R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����R��[
��U���7�2�;�u�w�}�W���Y�����D�����b�u�h�}�8�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V ��]���6�;�!�9�0�>�G������R��G�����4�
�:�&��2����Y�Ƽ�9��a1��*���|�n�u�u�2�9��������9l�N�U���&�2�7�1�`�d�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4��4�(�������@��Q��A���-�!�:�1�>�;�(��&���F�U�����u�u�u�u�w�}�WϿ�&����Q�� ]�I���}�%�6�;�#�1����H����C9��P1������&�`�3�:�i�W���Y������C�����3�
�c�
�e�`��������_��G��N���u�0�1�%�8�8��Զs���K��G1�����1�m�u�&�>�3�������KǻN�����2�7�1�m��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�
��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����R�
N�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u���(���	����O��N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�d�3�8�g�<����Y����V��C�U���4�
�<�
�$�,�$���¹��^9��V�����'�6�o�%�8�8�ǿ�&����Q��\��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��G���!�0�u�u�w�}�W���YӇ��@��T��*���&�d�3�8�g�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����0�
��&�f�;���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϿ�&����P��h=�����3�8�d�4�$�:�W�������K��N�����<�
�&�$���݁�
����R��P �����o�%�:�0�$�<�(���&����U��=N��U���<�_�u�u�w�}����	����l��h_�\ʡ�0�u�u�u�w�}�W�������T9��R��!���g�3�8�d�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�g�1�0�F��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��F���8�g�4�&�0�}����
���l�N��*���
�&�$���)�(���&����@��h����%�:�0�&�6���������OǻN�����_�u�u�u�w�;�_���
����W��X�����u�u�u�u�w�}�WϿ�&����P��h=�����3�8�g�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�f�3�:�o�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<�(���&����l5��D�����f�4�&�2�w�/����W���F�V�����&�$��
�#�����&����T��E��Oʥ�:�0�&�4��4�(���&����9F����ߊu�u�u�u�1�u��������lW��N�����u�u�u�u�w�}��������V��c1��A���8�f�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӇ��@��T��*���&�a�3�8�d�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����
����g9��1����4�&�2�u�%�>���T���F��h��*���$��
�!��.�(ہ�
����l��TN����0�&�4�
�>�����N��ƹF��R	�����u�u�u�3��-��������^�C��U���u�u�u�u�w�<�(���&����l5��D�����a�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������T9��R��!���`�3�8�a�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��Q��@ʴ�&�2�u�'�4�.�Y��s���R��^	������
�!�
�$��(�������A	��N�����&�4�
�<��9�(��P�����^ ךU���u�u�3�}�'�.��������F��R ��U���u�u�u�u�6�����
����g9��1�����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϿ�&����P��h=�����3�8�`�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���4�'�9�
�8�����Hʹ��V9��1��*��
�d�i�u�#�����&����\��R�� �&�2�0�}�%���������C9��h^��*ڊ� �m�a�%�~�n�^��Y����A��C1�����:�
�l�e�2�m����@ǹ��Z�B"��&����!��7�%�>�(�������
9��]����!�u�|�_�w�}��������l*��G1�*ڊ�
�
� �l�o�-�W��
����\��h����� �&�2�0��/�(���?����\	��W��*���
�
� �l�c�-�^�������]��G1��؊�e�3�
�m��n�^�ԜY�ƭ�A9��h(��*���%�d�
�
���(���@�ד� F�d��U���u�6�
����%�������V9��E��G��"�0�u�&�;�)�݁�&����V��^��H��r�u�9�0�]�}�W���Y����_��X�����d�
�
�
��(�N���	��ƹF��E�����'��:�
�n�o����K����
T��G]��H�ߊu�u�u�u�%���������C9��h^��*ڊ�
� �l�a�'�}����Q����G��^1����m�}�|�h�p�z�W������F�N��*������0�:�i�(���&����W��=N��U���
�!��'��2�(���K����lU��B1�@���u�h�_�u�w�}�W���0����r4��R��Aފ�
�
�0�
�f�}����Q����G��h�����e�d�e�u�w�l�^ϻ�
��ƹF�N�����!��'��8��N����֓�l ��\����u�u�4�'�;���������
9��R1��@���
�a�
�f�k�}�W���Y����A��C1�����:�
�l�e�2�m�E���&����CW��_��]���
�8�g�<�%�:�F��Q���A��N�����u�u�u�u�6�/��������\��1�����c�'�2�g�n�W�W�������l ��h"����
�
�
�
�"�d�C���Y���F�N���������2�0�Cف�&ù��T9��N�����&�9�!�%�>�/���A����[�I�����u�u�u�u�w�<����&����	��h_��E���e�g�3�
�g��F�ԜY�ƭ�A9��h(��*���%�d�
�
���(���@�ߓ� F�d��U���u�4�'�9��2�(���	����9��1��*��
�g�"�0�w�.����	����A��^�]���h�r�r�u�;�8�}���Y���R��[�����:�%�d�
���(���&����9F���*����'��:��d�E���H�ԓ�F9��1��U��_�u�u�u�w�/�(���?����\	��W��*���
� �l�m�'�}����Q����G��^1����m�}�|�h�p�z�W������F�N��*������0�:�i�(���&����S��=N��U���
�!��'��2�(���K����lU��B1�F���u�h�_�u�w�}�W���0����r4��R��Aފ�
�
�0�
�b�}����Q����G��h�����e�d�e�u�w�l�^ϻ�
��ƹF�N�����!��'��8��N����ד�l ��[����u�u�4�'�;���������
9��R1��A���
�b�
�f�k�}�W���Y����_9��s+��'���'�
�c�0�f�/���Aӑ��]F��R�����
�0�
�e�d�m�W���H����_��=N��U���u�'�
�!��/�;���&�ߓ�l��h��L���%�n�u�u�6�/��������\��1�����`�3�
�b��n�K���Y���F��[1��1����!�'�
�a�8�F���������YN�����8�g�<�'�0�l�N���P���A�R��U���u�u�u�4�%�1�(���&����lW��1��D���3�
�b�
�d�W�W�������VR��S�����
�
�
� �c�e����D�ο�T��C1����`�4�1�;� �4����&���� S��G�U���7�8�'�0�>�;�(��&���F��R	�����:�
�
� �o�l����Ӗ��
9��Z�����
�:�
�
�"�e�D���P���F��Z�����<�3�
�m��o�K�������T��C1��*��
�f�:�u��2�(���&����V��G�U���7�8�'�0�>�4����&����CT�
N�����3�:�
� �b�d����Ӊ��A ��@1��*��
�g�n�u�w�?��������l��h�� ��b�%�u�h���N�������]9��^1��*��
�g�4�1�9�:��������l ��Z�����_�u�u�4�%��(���A�ғ�F�F����
�0�
�d�o�<�Ϫ�	����Z9��hY�*��n�u�u�6�%�$����Mʹ��Z���*���'�2�d�e�w�3�W���&Ź��U��]��G��u�u�1�9�#�9����
�ד�F9��1��U��_�u�u�u�w�<��������]��1����g�u�=�;��<����&����R��F�U���d�|�0�&�w�}�W���YӴ��T��V�����&�'�2�d�d�f�W�������V��R��*���a�`�%�u�j�u��������T9��N��ʻ�!�6�'�,�>�;�(��&���9F������1�<�3�
�a��E��Y���D��F��*����'��:������A���R��X ��*���
�|�0�&�w�m�L���YӀ��l
��q��9���
�c��3��d�(��E��ƹF�N�����:�0�!�'������!����P��D1����`�u�=�;��8�(���K����F9�� 1��]���h�r�r�u�;�8�}���Y���\��h�����&�2�
� �a�l���Y����K��X
�����
�f��3��i�(��E��ƹF�N��*���g�`�8�-�>�;�(��&����[�������:�
�:�
��(�B���	����[�I�����u�u�u�u�w�-�!���&ƹ��U��^��F�ߠu�u�x�u�%��(߁�&����lT��h�����&�<�;�%�8�8����T�����h��*���
� �g�f�6�����
����C��T�����&�}�%�6�{�<�(���&����l5��D�����g�u�%�&�0�>����-����l ��h]��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y�έ�l��D�����
�u�u�%�$�:����&����GU��D��\ʺ�u�4�
�:�$�����&���R��^	������
�!�
�$��^���Y����l�N��U���u�2�%�3�g�;�D���&����R��RN�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�0�-�����Փ�F9��1��*���i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9l�N�����e�3�f�3��d�(���
����Z�P�����3�f�3�
�n���������C9��V�����_�u�u�'���(���&����
U��Y1�����d��i�u��<�E�������R��=N��U���
�
�
�
��(�E�������G��h8��Hʳ�%�;�1�
�2�0�B܁�&����V��d��Uʲ�%�3�e�3�d�;�(��&����R��h8��Hʥ�d�8�-��>����s���K��E�� ��e�%�u�&�>�3�������KǻN����� �f�e�%��.����	����	F��X��´�
�<�
�&�&��(���&����J��G1�����0�
��&�e�;���Y����Z��D��&���!�
�&�
�{��E�������G9��h]�*��u��
�
�����O����)��h8�� ��e�%�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N�����
�e�
�e�k�}�'݁�&����V��F�U���u�:�;�:�g�f�W���Y����_��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�d�|�#�8�W���Y���F�	��*���f�e�%�u�j��F���H����F9��1��]��x�d�1�"�#�}�^�ԜY���F��D��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}����s���F�N�����3�
�e�
�g�a�W���&����P��h��F���%�}�a�x�f�9� ���Y����F�N�����u�u�u�u�w�}�WϹ�	���� V��G^��H���������/���!����k>��o6��-���w�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����V��N�����u�'�6�&�y�p�}���Y����U��^��D���&�2�
�'�4�g��������C9��P1������&�d�3�:�m�W���
����@��d:��؊�&�
�y��f�����H������D�����
��&�`�1�0�C�ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��G1�����0�
��&�b�;���PӒ��]FǻN��U���u�u�'�
�"�n�G���Y����cW��h��*��e�f�u�u�w�2����I��ƹF�N�����u�}�%�6�9�)���������D�����
��&�g�1�0�F�������9F�N��U���u�'�
� �d�m����DӇ��P	��C1��Cފ�`�`�`�a�d�}�W�������V�=N��U���u�9�<�u��-��������Z��S�����2�6�0�
��.�F��������YNךU���u�u�u�u�%����I����[��G1�����9�c�
�f��h�_��T����\��XN�N���u�u�u�0�$�}�W���Y���F��E�� ��e�%�u�h�u��/���!����k>��o6��-�������u�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����U��^��G��u�!�
�:�>�����۔��Z��B �����}�!�
�:�>�����ە��]��P�����e�
�e�u�w�4����^���T��Q��Eڊ�d�|�y�c�~�f�W�������F9��1��U��2�%�3�
�g��E��Y����G	�G�U���<�
�<��%�����H����P��G\��Hʦ�1�9�2�6�!�>��������V��{1��*���
�:�%�<�%�:�E��Y�ƹ�@��R
�����;�!�9�g�f�t�}���Y����@��Q��G܊�g�i�u�&�0�?��������V��V �����c�
�
� �o�m����s���]��D�����<�3�
�a��o�K���	����Z9��h��M���%�u�'�&�0�?��������F9��1��\�ߊu�u�0�&�0�?����&����CU�
N��#���
�
� �a�g�-�_������\F��UךU���:�
�4�'�����@����[�Y�����<�
� �a�b�-�W���	����F
��1�����3�
�`�
�e�f�W�������A��h�����3�
�m�
�d�a�W���Y��� ��h �����'�
��4�4��(�������A��^�U���;�}�0�
�:��(���O�ӓ�N��S��D���0�&�u�u�w�}�Wϸ�	����V9��E��#���6��
�'�!��(���&����l�N�����:�
�
� �a�o����D�θ�C9��h��*��`�4�1�!�'�l�(�������V�=N��U���'�9�"�3��d�(��E����A��P��*��� �a�c�%�w�3�W���&����l ��Y�����_�u�u�x�w��(���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��v1�����9�
�;�&�0�<����&����\��E�����
�
�
�
�'�+����&ù��e9��h��*���2�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����8����C9��SG�����u�u�u�u�w�}�WϮ�I����l��A�����<�u�h�%�g��!���&����9F�N��U���0�_�u�u�w�}�W���&ù��e9��h��*���&�2�i�u���(���	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
���(���
����@��YN�����&�u�x�u�w�-�G���/����@��V�����'�6�o�%�8�8�Ǯ�I����F��1��#���0�y�%�e��������ƹF��R	�����u�u�u�3��<�(���
����T��N�������4�
�;�t�W������F�N��Uʥ�e���<��4�W��	�֓�l0��N��U���0�&�u�u�w�}�W���YӖ��l'��h�����i�u�
�
������s���F�R ����_�u�u�;�w�/����B���F��[�����'�i�u��9�9�(�������R��o>�����
�
�0�
�g�h�}���Y���C9��h=�����4�
�9�u�$�4�Ϯ�����F�=N��U���`��6�:��-��������]9��X��U���6�&�}�%�4�q��������V��c1��@���8�a�u�-�#�2�������� 9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����:�}�0�<�4�3�(�������l��
N��*���&�
�#�
�~�t�W������F�N��Uʥ�d�
�0�!�%�<�(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʥ�d�
�0�!�%�<�(���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&¹��K9��V�����;�&�2�4�$�:�W�������K��N�����8�-��4��1�(���
����@��Y1�����u�'�6�&���(���&����l��N��D���-��4�
�;�����s���Q��Yd��U���u�<�u�}�'�>��������lW���*���
�
�%�#�3�t����Y���F�N��U���
�4�
�
�'�+����&����[��h_�����
�%�#�1�]�}�W���Y����l�N��U���u�%�d�8�/���������l��R�����8�-��4��1�(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����8�-��<��4�W�������A	��D�X�ߊu�u�
�
�6��(���
����@��Y1�����u�'�6�&���(���&����lW��V��*���2�u�
�
�6��(������F�U�����u�u�u�<�w�u��������\��h_��U���
�4�
�
�'�+��������9F�N��U���u�
�
�4���������C9��Z��#�ߊu�u�u�u�;�8�}���Y���F�G1������<�
�<�w�`��������l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��8��������W9��h��U���<�;�%�:�2�.�W��Y����lT��R�����
�9�
�;�$�:��������\������}�
�
�0�>�9��������lT��R�����
�9�
�'�0�W�W�������F�N�����}�%�6�;�#�1����H����lT��R�����
�9�|�u�?�3�}���Y���F�G1��%���:�
�%�#�3�4�(���Y����lT��R�����
�9�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�0�<�3�<�(���&����Z�
N��G���'�:�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*؊�0�<�1�<��4�W�������A	��D�X�ߊu�u�
�
�2�4����&����R��P �����o�%�:�0�$�-�E���������h>�����%�0�y�%�e�����&����_�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�0�>�9�������G��d��U���u�u�u�%�e�����&����Z�
N��G���'�:�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�0�<�3�4�(���Y����lT��R�����0�n�u�u�w�}�������F�R �����0�&�_�u�w�-�Dׁ�&�ד�F9��1��U��}�4�'�
��(�O���	�ƭ�WF��Y	��*���
�;�&�g�%�:�F��P���F��V��*��� �a�`�%�w�`�_�������lR��h����&�2�7�!�%�:�N��B�����1�����4�
�
�
�"�e�F���Y���W��C�����&�d�3�
�g��Dϱ�Y����Q��1����e�|�_�u�w��N�������]9��Y�����
�`�
�g�k�}���&����A��h��*���m�d�%�u�8�}��������EW��UךU���
�
�
�<�>�:���E�ƭ�A9��h(��*���%�d�
�
���(���&����9l�N�U���
�
�<�<�0�8�G���&����R��P �����&�{�x�_�w�}�(ہ�&����]��h^�����1�4�&�2��/���	����@��G1��Yʴ�
�<�
�&�&��(���&����J��O�����<�3�
�c��o�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ�ӈ��N��^�����
� �c�f�'�}�W�������l
��h^��\���=�;�_�u�w�}�W���Y����f9��Z��*���
�%�#�1�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����h;�����2�0�e�4��1�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u���(�������lW�
N�����
�:�
�:�'�l�(݁�&¹��T9��UװU���x�u�
�
��4�����ד�C9��SN�����u�'�6�&�y�p�}���Y����f9��Z��*���
�%�#�1�6�.���������T��]���6�y�4�
�>�����*����9��Z1�U���!�:�1�<�1��A܁�K���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�(���&����]��X�����6�;�
�
�"�k�D���Y�ƭ�l��D��ۊ�|�|�u�=�9�W�W���Y���F��1��!���;�
�
�
�'�+���Y����\��h�����n�u�u�u�w�8����Y���F�N��*ފ�
�<�<�2�2�l���������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����q9��V�����;�&�2�4�$�:�W�������K��N�������4�
�;���������Z��G��U���'�6�&�}���(���	����F��1��#���
�9�
�'�0�W�W�������F�N�����}�%�6�;�#�1����H����lS��h8�����1�|�!�0�w�}�W���Y�����h,��*���#�1�<�
�>�}�JϮ�L����l��A�����u�u�u�9�2�W�W���Y���F��1��#���
�9�
�;�$�:�K���&ƹ��e9��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����Z��^	�����;�%�:�0�$�}�Z���YӖ��l$��h�����4�&�2�
�%�>�MϮ�������h,��Yʥ�`���%�2�q����;����C9��SGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�`���������G��d��U���u�u�u�%�b��!���&����[��h[��*��u�u�u�u�2�.�W���Y���F���*���
�;�&�2�k�}�(ځ�&����V��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʥ�c���8�9��(���DӅ��z(��o/�����
�a�0�e�%�:�E��s���K�G1��#���8�;�
�
��-��������]F��X�����x�u�u�%�a��#�������9��h��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�h����M�Ʃ�Z��Y
��*���c�f�%�|�w�}�������F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���`�3�8�a�w�3�W���Qۃ��G��S1�����c�
�g�h�6�����&����O�N�����u�u�u�u�w�}����/����Z��R1�����9�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����e9��Z��*���
�%�#�1�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R�����u�%�c���0����&�����~ ��-���!�'�
�a�2�l����K����9F�C������8�;���(�������@��YN�����&�u�x�u�w�-�A���-����T9��1��*���
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	��������F��^�����
� �c�f�'�t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�`�3�:�i�W���Y������C�����3�
�c�
�e�`��������_��G��\ʡ�0�u�u�u�w�}�W���	�Г�l2��^ �����4�
�9�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���C9��a1�����
�
�
�%�!�9�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�@���/����E
��^ �����&�<�;�%�8�8����T�����h-��*���#�1�<�
�>���������PF��G�����%�b���6����	�ѓ�l0��G1�����0�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���&����R��[
��U���;�_�u�u�w�}�W���&Ĺ��e9��h��*���&�2�i�u���(���	����l�N��Uʰ�&�u�u�u�w�}�W���	�ѓ�l0��G1�����
�<�u�h�'�j�4�������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�`��!���&����R��P �����&�{�x�_�w�}�(؁�&����l��h�����%�:�u�u�%�>����&Ĺ��eJ��hY��*���'�2�u�
���(������F�U�����u�u�u�<�w�u��������\��h_��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�
�9�.���Y����p9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��a1��*���u�h�%�b������B���F���U���u�u�u�0�3�-����
��ƹF��hV��*���<�2�0�e�k�}����=����a��Z1�*���
�0�
�e�l�W�W���TӖ��l1��^�����e�4�
�9�w�.����	����@�CךU���
�
�
�<�>�:��������W9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�
�&��q��������Z9��hX�*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C[�����|�4�1�;�#�u��������l ��X�����u�%�6�;�#�1�F��P����[��=N��U���u�u�u�
����������l��A��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�-�O�������T9��1��*���u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǻN��*Ҋ�
�<�<�2�2�l�K�������v>��e����
�
�
�0��k�L�ԜY�����h9�����2�0�d�4��1�W�������A	��D�X�ߊu�u�
�
��4�����ד�C9��S1�����
�'�6�o�'�2��������F��h��*���$��
�!��.�(������\��^1��*��
�g�_�u�w�8��ԜY���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��ߊ�&�
�|�4�3�3��������]��h��C���%�u�u�%�4�3����H���O��_�����u�u�u�u�w��(�������l��h�����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϮ�A����Z��P1��D���
�9�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���
�0� �!�e��(���N�ӓ�F�	��*���f�e�%�}�d�9� ���Y���9F������!�f�<�;�#�;�(��&���F��Z��B���2�d�e�u�8�}��������EW��UךU���
�4�g�g�e�0��������9��R�����u�u�u�
�6�o�Bց�����l��@��U·�8�'�0�<�>�3��������9��^��H��r�u�9�0�]�}�W���Y����\��h��G������n�w�}��������l ��\�����h�&�1�9�0�>�����ο�Z ��[��]���<�;�1�%�g��!���&������^ ����� �&�2�0��m�W���	����@��A]��D��x�u�:�;�8�m�^���B�����V��@ފ� �`�e�%�w�`��������9��X����!�u�g�n�w�}��������l ��_�����h�&�1�9�0�>�����ι�@��R
��*���g�`�
� �b�m����Rӓ��Z��SF����
�
� �c�o�-�^��Y����l0��1�*���b�`�%�u�j�.��������V��EF�����0�}�
�4�e�h�(���&����F�B �����}�8�
�l�>�;�(��&���l�N��#���
�
�
� �b�m����D���F�N��*���&�
�#�g�o�m�G��Y����N��S�����3�
�e�
�e�m�W���H����_��=N��U���u�
�4�g�`�;�(��&����F�G1��؊�
� �
�
�"�h�E���Y���F�N�����:�&�
�#�e�j�1���?�ƻ�V�U�����<�<�<�3��l�(��I���W����ߊu�u�u�u��<�E�������9��d��Uʥ��9�
�e�1��Oށ�J���9F�N��U���4�g�g�g�:�%����&����CU��_��]���0�2�
�
�"�e�N���Q���A��N�����u�u�u�u�'��݁�&����U��UךU���
�4�g�c�1��C؁�H���T��Q��Eڊ�g�c�u�u�w�2����I��ƹF��h8��G���3�
�f�
�e�a�W���&����P9��T��]���<�;�1�%��1�(ف�����R�N�����0�}�8�
�����N����]ǻN��*���g�<�3�
�`��D��Y���F������!�9�f�
�w�5��������P9��hV�*��e�u�u�d�~�8����Y���F��h8��G���
� �b�`�'�f�W���	����9��Q��F܊�f�i�u�u�w�}�WϿ�&����G9��\��3�����"�0�w�2��������U��\��G��u�u�d�|�2�.�W���Y�����V��@ߊ�0�
�e�e�]�}�W�������Z9��hZ�*��i�u�1�9�#�9����
����P��G\�����%�6�;�!�;�l�F��Y����Q9��D��*ފ� �f�b�%�w�`�_���&����U��_��Gʴ�1�$�<�
�"�n�@���P���F��h�����c�3�
�e��o�K�������9��Q��L܊�g�4�1�$�>��(���L�֓� O��N�����&�<�;�m�1��@؁�K�����h��M���2�d�g�u�9�}����J����lW��G�U���$�<�
�
�"�h�G���Y����A��B1�E���}�d�1�"�#�}�F��Y����Q��Q��@݊�d�i�u�'��(�D���	����K�
�����e�n�u�u�&�4�(���J�ѓ� F������
�`�
�d�e�}��������l�N��G���
�m�
�g�k�}�G������G�� _�� ���m�%�u�u�'�>��������O��[��W���_�u�u�
��(�@���	���D�������8�
�c�3��o�(��DӇ��P	��C1��G݊�|�0�&�u�f�f�W�������l ��^�����h�&�1�9�0�>�����ο�T����*ߊ�
� �a�f�'�t�Zϭ�����G��^1��*��
�d�|�_�w�}�(���&����W��N�U���
�:�<�
�2�)�ǭ�����G�� 1�����d�
�d�u�w�4��������l��B1�B���|�n�u�u�%�����K����Z�D�����6�#�6�:��4��������l ��_�����x�&�2�0��0�(ށ�&����^��G����u�
� �f�n�-�W��[����[����*���3�
�c�
�f�`��������_��h^�����u�d�n�u�w�/����&����lS��h�I���!�%�b�
�"�h�O���Y����lT��B1�G���|�_�u�u���(�������
9��R��]���
�m�3�
�c��Dϱ�Y����U��Y��G��u�u�'�<�>�4����@¹��Z���*���3�
�m�
�d�2�W�������l��d��Uʦ�9�!�%�
��(�A���	���D��������9�
�:��2��������W������!�9�g�e�w�1����[���F��[1�����3�
�b�
�e�a�W��Y����N��h��3����:�
�
�2��O���Y����\��h��*���0�&�u�e�l�}�Wϭ�����l ��]�����h�2�%�3��m�(��O���F��@ ��U���_�u�u�<�9�4�(���&����l^��h�I���&�2�7�!�e�/���I�ƴ�AF��h�����#�
�|�_�w�}���&����V��N�U»�"�<�;�<��(�C���	�ƣ���h��F���
�b�
�g�l�}�WϪ�	����Z9��hX�*��i�u�!�
�8�4�(�������V��RF�����0�}�7�4�$�:�(ف�����l��]�\�ߊu�u�8�
�e�4����KŹ��Z�	��*���f�c�%�u�8�}��������EW��UךU���u�u�8�
�����A����[��C
�����
�0�!�'�%�.����������h-��*���&�2�y�f�~�W�W�������l��B1�B���u�h�&�1�;�:��������A��M�����;�1�$�
�$�4��������W��]�\�ߊu�u�8�
�n�4����A¹��Z�D�����6�#�6�:��8��������]��F�����;�m�3�
�`��E��K����F�N�����`�<�3�
�g��F��Y����_	��T1�����}�0�<�0�$�:����&����lS��Q��GҊ�g�y�f�|�]�}�WϪ�	����Z9��hY�*��i�u�!�%�`����I����K	��V�����
�#�
�|�]�}�W���&�ד�l ��\�����h�}�
�m�>�4�(���A�ӓ�F��EN��*���&�
�#�
�~�W�W�������l ��X�����h�2�%�3��m�(��O���F��@ ��U���_�u�u�8��k����Oƹ��Z�C��C܊� �f�`�%��j�Z������\F��d��Uʡ�%�c�
� �d�h����DӁ��l ��^�����d�x�d�1� �)�W���s���G��V�� ��f�%�u�h�0�-����Iù��P��N����!�u�|�_�w�}����A���� ^��G]��Hʡ�%�c�
� �d�n����Aӂ��]��V����u�8�
�
��(�C���	���N��@�����
� �a�`�'�}����	����@��A_��\�ߊu�u�8�
�f�;�(��&���F��G1��*��
�g�f�u�w�}�������9F���*���3�
�m�
�d�a�W���&����V��F�U���;�:�f�|�]�}�W���&�Г�F9��1��U��2�%�3�
�g��E��Y����W	��C��\�ߊu�u�8�
�o�;�(��&���F��G1��*��
�g�g�u�8�3���P���F��G1�*���b�e�%�u�j�-�!���&�ߓ�F9��1��]��1�"�!�u�f�f�W���Y����^��h�� ��f�%�u�h�$�9��������G	��E�����<�;�1�'��n����IĹ��J��G����u�u�u�8���(���M�ѓ�F���*���<�
�0�!�%�/����Q����V��hY��*���;�&�2�y�c�t�}���YӒ��l��X�����
�e�
�g�k�}���&����U�� [��Gʺ�u�'�0�2�c���������l��B1�M���|�_�u�u�:��(�������9��R��]���;�<�
�0��d�W���Y����\��h��*���_�u�u�u�w�0�(�������l��S�����:�<�
�0�#�/�����ο�T����*���
�;�&�2�{�n�^�ԶY����9��b,�� ��� �!�4�!�d����@����[��C
�����
�0�!�'�"�.����Q����c��X
�����2�u�u�;�>�3�Ǯ�/����V��B1�D���|�n�u�u�"�9��������V��G\��H���8�
�0�:�0�3����I�����������
�0�
�l�~�W�W�������_	��Y�����
�g�
�g�k�}����I����T��G\��ʥ�f�
�
�
�"�i�B���P���WF��_��