-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�_�&�w�8��������Z��X����_�0�!�!�w��B���8����l��X��C޻�
�g�g�<�]�}�W�������l�N��Uʜ�u�u�u�u�w�}��������W��=N��U���u� �
���}�MϷ�����\�UךU���u�u�<�e� ��?������V�
N�N���u�u�u�1�"��>���Y�ƥ�G��EN�U��u�u�|�_�w�}����Q���F���U���u�;�u�!��2���Y���F��R��U���;�u�!�
�8�4�L���Y�����N��U���u�!�
�:�>�f�W���Y����Z��T�����!�
�:�<��8��������d/��C����!�u�|�_�w�}�W������	F��CN�����2�6�#�6�8�u����.����W��X����_�u�u�n�2�9������ƓR��^�����u�'�=�:�w��B���8����l��X��C޻�
�g�g�<�]�}�W��T���K�C�X���x��8�:�2�)�Z��T���K�C�X���_�u�u�:�'�3����<�Ӎ�v'��h^�����!�3�
�
�8�9���Y��ƹF�N�����}�u�u�u�w�}�Wϭ�����R9��V��U���u�o�<�u�$�9�������F�N��Uʦ�4�<�
�
�3�)�W���Y����Z�D�����6�#�6�:��n��������l�N��U���u�8�4�<��8��������WF��X�����9�2�6�_�w�}�W���Y�ơ�R��h�� ���!�4�4�u�w�(�W���&����P9��T��]��1�"�!�u�~�}�W���Y����F�R �����:�0�!�_�w�}�Z��T���K�C�X����6�9�&�0�<�W��T���K�C�X�ߊu�u�<�;�;�<���������h����u�u�&�2�6�}�(������	F��S1�����#�6�:�}�d�9� ���Y����F�D�����
�#�9�1�w�}��������9F������'�!�4�4�w�g��������l��C��F���:�;�:�e�l�}�Wϭ�����W��h��D��&�1�9�2�4�+����Q����l1��c&��U���;�:�e�n�5�:����Y���K�C�X���x�x�x�u�9�)��������K�C�X���x�x�x�u�w�0�Gڟ�<����9��h�����e�;�
�&��i�������]����@����3�e�4��4����I����W��ZךU���:�!�8�%��}�W���Yӕ��K��V1�����u�u�u�h�w��������F�N�����
�
�1�!�w�}�W���GӇ��W��d��U���u�8�4�<��8��������WF������1�_�u�u�w�}�(���
����F
��C
�����k�'�!�4�6�}�W���s���K�C�X���x�x�x�x�z�}��������K�C�X���x�x�x�x�z�}�WϿ�����WF�I�N���u�4�!�4�6�}�J����֓�z"��_�����:�e�h�u�g�t� ���Y�Ψ�]V��B�H���1�;�
���p�W������[�6��\���'�}�<�e�5�;�W���Y����l1��c&��U���;�:�e�h�w��^�������W��h��D�ߊu�u�:�!�w�}�K���&����R]ǑN��X���x�x�x�x�z�p�Z��Tӯ��F��B�����x�x�x�x�z�p�Z��s���C��R��]���|�7�2�;�w�}�W����Ư�XA��R �����6�>�h�r�p�)��ԜY���F�N��U���h�r�r�!�2�W�W���Y���F�N��ڊ� �d�i�u�>�m�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�;�u�'�?�)������