-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�_�&�w�8��������Z��X����_�0�!�!�w��B���8����l ��S����;�
�g�&�d��(���������N�����'�6�}�u�w�}�Wϗ�Y���F�N�����'�o�u�n�w�}�W���7����g'��N����2�'�o�u�l�}�W���Yӂ��9��s:��Oʼ�!�2�'�o�w�o�}���Y���W��h9��!���u�;�0�0�w�`�D��Y���F��X��"����o�<�!�0�/�M���K���O��N�����u�_�u�u�w�}����Y����]F��C
�����n�u�u�u�w�/����Y�ƥ�F��S1�����_�u�u�u�w�8�W���Cӏ����h����u�u�u�u�3�3�W���Y���@��[�����6�:�}�<�g�
�3���Hӂ��]��G�U���u�u�1�;�w�}�W���Y����_	��T1�����}�<�d����FϺ�����O��N��U���:�6�1�u�w�3�W���&����P9��T��]���:�;�:�e�l�}�W���Yӂ��GF�N��ʦ�1�9�2�6�!�>��������z"��_�����:�e�_�u�w�f��������J]ǑV�����!�'�u�'�?�2�W���L�щ�p ��h�����7�f�;�
�e�.�D݁�&����l����U���x�x�x�x�z�p�Z��T���%��G�����x�x�x�x�z�p�Z��T���F�T�����!�8�e����(߁�	����W ��U1�����
�&�
�g�>�W�W���Y�Ƽ�A�=N��U���u�u�u�6�<�}�W���Y���F�N��Oʼ�u�&�1�9�0�>�}���Y���F�V�����u�u�u�u�w�}�W���Cӏ����h����u�u�u�u�w�}��������G��^
��U���u�u�u�;�w�)�(�����ƹF�N��U���
�-�&�4�#�<����Y���F��^ �����9�2�6�#�4�2�_������\F��d��U���u�u�u�&�6�4�(�������F�N��U���;�u�!�
�8�4�L���Y���F������7�!�4�4�w�}�W���Y�ƥ�F��S1�����#�6�:�}�f�9� ���Y����F�N��U���&�4�<�
�'�/����&����Z���U���
�:�<�n�w�}�W���Y����l��D1�����<�;�!�4�6�}�W���Y����_	��T1�����}�u�:�;�8�m�L���Y���F������'�&�9�
�!�1����Y�ƣ�GF��S1�����_�u�u�u�w�}�W�������V��C1�����u�u�o�:�#�.��������V��EF�U���;�:�e�_�w�}�W���B����������;�n�u�u�z�p�Z��T���K�C�U���4�u�<�;�;�p�Z��T���K�C�U���&�2�4�u�4�6�W���Y����@��[���ߊu�u�<�;�;�<����Y���\��C
�����n�u�u�&�0�<�W�������F�N�����2�6�_�u�w�4��������G�N��U���
�:�<�
�2�)���Y����G	�UךU���<�;�9�7�#�<����Y����G��X	��N���u�&�2�4�w�����Y���	F��S1�����#�6�:�}�f�9� ���Y����F�D�����%�!�4�<�w�}�W���&����P]ǻN�����9�:�
�1�#�}�W��
����\��h�����b�1�"�!�w�t�}���Y����R
��h�����u�u�u�!��2���Y����Z��[N�����4�u�u�o�$�9��������G	��_�����:�e�n�u�w�.����Y����l��N��Oʦ�1�9�2�6�!�>�����֓�z"��_�����:�e�n�u�w�.����Y����l��N��Oʦ�1�9�2�6�!�>�����ד�z"��_�����:�e�n�u�w�.����Y����W��B�Oʦ�1�9�2�6�!�>����Y����G	�U�����_�u�u�x�z�p�Z��T���K�N�����!�4�<�;�z�p�Z��T���K�=N��U���`�b��3�g�<�(�������lW��B�����f�
�u�u�8�-����Y����rQ��t��*���3�1�3� ����������l�N�����4�u�_�u�w�}�W������F�N��U���u�u�h�u�4�6�}���Y���R��R ��U���u�u�u�u�w�}�J�������l�N��Uʦ�4�<�
�
�!�1����Y���[�V1�����y�u�u�u�w�.����&����R��N��U���u�k�4�!�6�<�}���Y���@9��^��*���9�1�u�u�w�}�J���&����Z�N��U���&�4�<�
��9����Y���F�	N�����4�_�u�u�w�}�(���
����A��X �����1�h�u�%�#�<���Y���F��h�����0�4�<�;�#�<����GӉ��G��VBךU���u�u�
�-�$�/����&����Z�N��U���#�9�1�_�w�}�W���&����l��B�����4�u�u�h�w�����s���]ǑN��X���x�x�x�x�z�p�Z��Tӧ��Z��R ��X���x�x�x�x�z�p�Z��s���R��N��U��u�9�n�u�w�<����Y���F��d��Uʴ�!�4�<�u�k�}�F��Y����l��C��U��}�<�e����FϺ�����F�I�\ʢ�0�u�}�<�g�?����Y�ƨ�]V��~*��X���:�;�:�e�j�}�/���YӉ����1�����u�u�<�e� ��?������\F��
P�� ���|�0�&�u�>�m����B�����A�����h�r�r�_�w�}�(������[�S��*����x�u�:�9�2�G��Y�����YN�����
� �d�h��9�ށ�0����F��@ ��U���k�r�r�|�w�/�_���H����F�N��ۊ���x�u�8�3���D����O���ʱ�;�
� �d�]�}�W�������WF�I�N���u�:�
�1�#�}�K���I����V�������:�6�1�
�"�l�J���!����AF��G�����3�u�u� �u�t����Y���V��L��U���:�0�7�3�~�W�W������F�S��*���!�n�_�u�w�p�Z��T���K�C�Xʜ�%�!�7�3�2�}�Z��T���K�C����u�'�6�&�w�>��������F�N�����9�r�#�;�w�3�W���Y���F��R ךU���u�u�u�u�1�>�W���H�Ƹ�VǻN��U���u�u�u�u�>�m����Y�����UךU���u�u�u�u�w�}��������F�
��D�ߊu�u�u�u�w�}�W���	����l��N�U���:�0�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=��U���=�!�6� �2�W