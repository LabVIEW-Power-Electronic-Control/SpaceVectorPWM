-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�m�m�d�a��}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e�4�%�4�m��W���&����p9��t:��U��u�:�;�:�g�f�W�������\��yN��1�����_�u�w��(�������l��T��;ʆ�����]�}�W���&����	F��=��*����
����u�FϺ�����O��N�����8�-�4�
�;�}�W���*����|!��d��Uʥ�g��'�:�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����c��X
�����1�o��u���8���B�����h;�����2�0�e�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���&ǹ��g��Y	��*ڊ�%�#�1�o��	�$���5����l�N��A����8�;�
��}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y����lR��h:�����0�d�4�
�;�}�W���Y����)��tUךU���
�
�0�4�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ӓ�V��V�����u������4�ԜY�Ƽ�9��c�����
�u�u� �w�	�(���0����p2��F�U���;�:�e�n�w�}����/����Z��R1�����9�u�u� �w�	�(���0��ƹF��hX��*���<�2�0�d�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����e9��Z��*���
�%�#�1�m��#ύ�=����z%��N������!�8�;���W���,�Ɵ�w9��p'��#����u�f�u�8�3���B�����h9�����2�0�e�4��1�W���,�Ɵ�w9��p'�����u�
�
�
�>�4����H����f2��c*��:���
�����l��������l�N��M���!�8�;�
����������f2��c*��:���n�u�u�%�f���������f2��c*��:���
�����}�������9F���@���6�:�
�%�!�9�Mϑ�-ӵ��l*��~-��N��1�_�_�'�?�)����ӄ��R��QN��M��d�a�
�u�$�W�W�������F��t!��*���������W���-����l�N����� �0�����2���0����} ��X�����u�u�'�=�#�>�������F��qV��Dۑ�3�e�=�&�>��G���Mߝ��`9��g;��!���h�-�y����"���5����J��d1��%������e���>���-����g[�� �E���a�a�d����'���:����T��^�E����
�� ���?ұ�����{*��d7��6����g�{�b�g�m�?���*����r2�B��&������;�9�q�;��� ����~[��"��&�����d�y���.���?����J��d1��;����m�`�(�l�}�WϽ�����GF��h�����:�<�
�u�w�	�(���0����A��d��Uʶ�;�!�;�u�'�>��������lV�=��*����u�h�r�p�W�W�������]��G1��*���
�&�
�u�w�	�(���0����p2��F����!�u�|�o�w�m�F��Y����\��V ������&�g�3�:�l�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���H����F�T�����u�%��
�#�����Y�Ɵ�w9��p'��#����u�g�1� �)�W���C���V�=N��U���&�4�!�4��2�����ԓ�\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����F��d:��9�������w�m��������\�_�����u�:�&�4�#�<�(���
���� T��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��h\��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�D���_�u�u�&�0�<�W���:����^F��d:��9�������w�o��������\�^�W�ߊu�u�!�'�5�)�W���&����W��T�����2�_�u�u�#�/����Y����V��S��U���4�
��3�:�g�����ƥ�D��Y�����u�<�;�9�6�����
����g9��1����o������}���Y����R
��G1�����1�d�u�u���6��Y����Z��[N��E���%�4�<�
�>�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�����%�0�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�u�W�W���������h�����%�#�1�<��4�W���-����t/��=N��U���;�9�%�e�6�-����&����C��T��!�����u�h�p�z�}���Y����R
��h_�����;�&�2�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��l��h����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�n�u�u�$�:����&¹��K9��h��*���&�2�o����0���s���@��V��*ۊ�4�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���&����\��Y1����������4���Y����W	��C��\�ߊu�u�<�;�;�-�E�������C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�<�;�;�-�E�������R��[
�����2�o�����4�ԜY�ƿ�T����*���<�1�4�
�;�����Cӵ��l*��~-��H��r�_�u�u�>�3�Ϯ�L����R9��h��U����
�����#���Q����\��XN�N���u�&�2�4�w��(�������TF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���&�2�4�u����������W9��h��U����
���l�}�Wϭ�����C9��U��*���#�1�%�0�w�}�#���6����	[�I�U���&�2�4�u�'�.��������	F��x"��;�ߊu�u�<�;�;�;�(�������^9��z/�����!���&�%�:�E��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����2�6�0�
��.�E������5��h"��<��u�u�&�2�6�}��������lW��T��:����n�u�u�$�:��������9��1��*��
�%�1�;�w�}�#���6����9F������3�
�:�0�#�/�(���8����q��d)�����'�2�g�`�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������`9��S�������9�=��)�$���
�ԓ�V��^��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u��3��������e+��G������
�
�0��n�W���-����t/��a+��:���b�1�"�!�w�t�}���Y����R
��E��*ڊ�
�
� �d�e�<�(�������`2��{!��6�ߊu�u�<�;�;�:����I����l ��]�����1�0�o����0���s���@��V�����
�
�
�
�"�l�E���&����JF��d:��9����_�u�u�>�3�Ϲ�	����l ��h��D���<�
�9�=��}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��E���d�3�
�f��3����K����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�
��(�F�������G��T��!�����
����_������\F��d��Uʦ�2�4�u�'���(���&���� T��G1�����
�u�u����>���<����N��
�����e�n�u�u�$�:��������9��1��*��
�%�'�!�%��W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����3�d�3�
�d���������F��d:��9�������w�n�W������]ǻN�����9�2�%�3�g�;�F���&����R��R����o������!���6�����Y��E��u�u�&�2�6�}����&ù��9��h_�*���6�u�u����>��Y����Z��[N�����e�3�g�3��i�(���
����\��c*��:���n�u�u�&�0�<�W���&����U9��Q��A؊�%�1�;�u�w�	�(���0��ƹF��^	��ʲ�%�3�e�3�e�;�(��&����W
��N��1�����_�u�w�4��������lV��h\�� ��g�4�
�0�3�}�W���&����p]ǻN�����9�2�%�3�g�;�E���&����Z��G�����e�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����l ��h��D���<�
�0�<�3�n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E��*ڊ�
�
� �d�e�4�(�������lW�=��*����
����u�FϺ�����O��N�����4�u�'�
���(݁�����l��`�����
�u�u����>���<����N��
�����e�n�u�u�$�:��������9��1��*��
�%�'�!�%��W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����3�g�3�
�c���������F��d:��9�������w�n�W������]ǻN�����9�2�%�3�g�;�E���&����R��R����o������!���6���F��@ ��U���_�u�u�<�9�1�����֓�lT��B1�G���
�0� �;�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��*���
� �d�g�6��������5��h"��<������}�f�9� ���Y����F�D�����'�
�
�
�����K����A��E ��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���&����U��\�����u�u��
���L���Yӕ��]��V�����&�$��
�#�����Y�Ɵ�w9��p'�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1�����֓�lW��B1�G���
�!�'�
�'�.�������5��h"��<���h�r�r�_�w�}����Ӂ��l ��h��*���d�g�4�
�#�/�(���
����l��T��!�����u�h�p�z�}���Y����R
��G1��*���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������W9��T��:����n�u�u�$�:����	����l��h_�U������n�w�}�����ƭ�l��h��*��o�����W�W���������D�����`�u�u����L���Yӕ��]��V�����1�
�m�o���2���s�����G�������d��1�m���0���F��E�����u�u�u�%�4�6�Mϗ�Y����)��tUךU���u�u�%�'�#�g�>���-����t/��=N��U���u�%�&�4�#�g�>���-����t/��=N��U���u�%�1�;�w�}�"���-����t/��=N��U���u�%�<�9�w�}�"���-����t/��=N��U���u�%�'�4�.�g�8���*����|!��d��U���u�<�
�9�?��W���7ӵ��l*��~-��0����}�d�1� �)�W���s���F�^ �����u�u�����0���/����aF�N�����u�|�_�u�w�}�W�������F��~ ��!�����
����_������\F��d��U���u�4�
�0�"�3�G��6����g"��x)��*�����}�d�3�*����P���F�N��*��� �;�d�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���Y�ƭ�l��B��G��������4���:����U��S�����|�_�u�u�w�}�������� F��x;��&���������W������\F��d��U���u�4�
�0�m��W���&����pF�=N��U���u�:�%�;�9�f�}���YӅ��C	��Y��3җ�d��3�e�1�o�>�ԜY�Ƽ�A�=N��U���u�%�6�>�m��W���&����p]ǻN��U���%�'�!�o��}�#���6����9F�N��U���&�4�!�o��}�#���6����9F�N��U���1�;�u�u��}�#���6����9F�N��U���<�9�u�u��}�#���6����9F�N��U���'�4�,�o��	�$���5����l�N��Uʼ�
�%�'�0�#�m�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y���F��Y1�����
�u�u����;���:����g)��]����!�u�|�_�w�}�W�������A��C1�Oʜ�u��
����2���+������Y��E��u�u�u�u�>���������\��yN��1��������}�D�������V�=N��U���u�%�'�!�%��W���,�Ɵ�w9��p'��#����u�f�u�8�3���B���F������'�
�u�u��}�#���6����e#��x<��F���:�;�:�e�l�}�W���YӇ��A��E ��U��� �u��
���(���-��� W��X����n�u�u�u�w�<�(�������\��b:��!�����
����_������\F��d��U���u�4�
�0�"�3�C��6����g"��x)��*�����}�d�3�*����P���F�N��*��� �;�`�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���Y�ƭ�l��N��U���
���u�l�}�Wϻ�Ӆ��C	��Y����0�<�_�u�w�/�(���&����U��\��U���%�;�;�u���Fޚ��֓�lWǻN�����8�%�}�u�w�}�WϿ�&����X��G1���ߊu�u�u�u�'�/���Y����@�N��U���4�
�!�'�w�c�����֓�lW��B1�G���
�!�'�y�w�}�W�������]�	N�����e�3�d�3��n�(�������9F�N��U���<�9�u�k�0�-�����ד�F9��1��*���0�_�u�u�w�}�������F��G1��E���d�3�
�f��-���� ���F�N��*���=�
�u�k�0�-�����ד�F9��1��*���=�
�y�u�w�}�WϷ�&����F�	��*���
�
�
� �f�o��������9F�N��U���7�!�
�u�i�:����I����l ��]�����0�4�e�_�w�}�W���	����F��N��U���
�
�
�
��(�F�������G��h^�U���u�u�4�
�2�(���D�ƫ�C9��1��D���
�f�
�%�%�)����U���F������'�
�u�k�0�-�����ד�F9��1��*��� �;�g�_�w�}�W���	����F��N��U���
�
�
�
��(�F�������G��h]�U���u�u�4�
�2�`�W���&����U9��Q��F؊�%�6�|�_�w�}�����֓�lT��B1�G��6�8�:�0�#�0�O��H�Ҫ�9��d��Uʥ�'�u�4�u�]�}�W���Y����_�	N��*���y�u�u�u�w�<�(���Y����C9��CBךU���u�u�%�&�6�)�J�������9��1��*��
�%�&�4�#�W�W���Y�ƭ�l��RN��U���
�
�
�
��(�F�������]�N��U���4�
�1�0�j�}����&ù��9��h_�*���<�9�y�u�w�}�WϿ�&����JF�	��*���
�
�
� �f�o��������9F�N��U��� �0�6�;��}�IϹ�	����l ��h��D���<�
�%�'�2�)�G�ԜY���F��h>�����f�h�u�'���(���&����T��Y1�����
�y�u�u�w�}����	����]��S����3�e�3�g�1��C݁�����A��C1����u�u�u�;� �8����&�����h��*���
� �d�g�>���������l�N��Uʴ�
�0� �;�g�`�W���&����U9��Q��A؊�%�'�!�'��q�W���Y����C9��C��*���k�2�%�3�g�;�E���&����R��R����_�u�u�u�w�-��������X��E��*ڊ�
�
� �d�e�<�(�������l�N��Uʴ�
�0� �;�d�`�W���&����U9��Q��A؊�%�'�!�'��q�W���Y����C9��C��*���k�2�%�3�g�;�E���&����R��R����_�u�u�u�w�-��������X��E��*ڊ�
�
� �d�e�<�(�������l�N��Uʴ�
�0�h�u�%��(߁�&����lW��h�����_�_�_�u�w�p�W���Y����V��D�����%��
�&�~�2�W���Y����VF��T�����x�u�u�4����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��G1��*���u�h�4�
��.�F�������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��=N��U���u�u�u�u�w�}�W���:����^F���;���&�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�P�����3�d�3�
�d���������C9��V�����4�&�2�u�%�>���T���F��G1��E���d�3�
�f��-��������@��C1�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�2�'�;�G���H����U��V�����
�%�&�4�#�/���Y����\��h�����n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}����PӇ���������7�1�l�|�~�)����Y���F�N��U���u�u�'�
���(ށ�����l��D�����
�!�'�
�2�}�JϿ�&����G9��P��D�ߊu�u�u�u�w�}�W�������N��h�����:�<�
�u�w�/�(���&����U��\�����4�,�|�!�2�}�W���Y���F�N��U���'�
�
�
�����K����@��C1��*���'�
�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W������lV��h\�� ��g�4�
�!�%���������V��D��ʥ�:�0�&�u�z�}�WϹ�	����l ��h��D���4�
�!�'��-��������l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�
�
�
��(�F�������R��V�����
�0�u�h�6�����&����P9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���g�3�8�d�w�3�W���Qۇ��P	��C1�����e�h�2�%�1�m��������9��h
�����|�!�0�u�w�}�W���Y���F�N�����
�
�
�
�"�l�E���&����G9��h�����0�u�h�4��2��������]ǻN��U���u�u�u�u�;�4�W���	����@��X	��*���u�'�
�
���(���H�ԓ�C9��V
��\ʡ�0�u�u�u�w�}�W���Y���F��E��*ڊ�
�
� �d�e�<�(�������l��E�����h�4�
�:�$�����&��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m��������E
��G��U���<�;�%�:�2�.�W��Y����lV��[��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����R
��V1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�0�$�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���Yӏ����D�����d�d�u�=�9�W�W���Y���F�N��U���u�%�e�4�'�<��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&���G��d��U���u�u�u�u�w�}�W���YӖ��l��_�����1�%�0�u�j�-�G���	����C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(߁�����C�������%�:�0�&�w�p�W���	�֓�_��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�g�<����	����[��G1�����9�f�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʥ�e�4�%�4�6���������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�~�)����Y���F�N��U���u�u�
�
�;�5�(������C9��V���ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lW��V�����1�%�0�u�$�4�Ϯ�����F�=N��U���
�4�
�%�!�9����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����2�7�1�d�f�}����s���F�N��U���u�u�u�u�'�l��������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&����P�C��U���u�u�u�u�w�}�W���Y�����h��*���#�1�%�0�w�`��������C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(ށ�����V��D��ʥ�:�0�&�u�z�}�WϮ�H����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�d�8�/�-����DӇ��P	��C1��F؊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����^��V�����|�!�0�u�w�}�W���Y���F�N��*ۊ�4�
�'�2�k�}�(ށ���ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�o�'�������l��h��ʴ�&�2�u�'�4�.�Y��s���C9��g�����%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��E��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z �V�����1�
�b�|�#�8�W���Y���F�N��U���u�u�u�
��8��������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&����S�C��U���u�u�u�u�w�}�W���Y�����h>�����4�
�9�
�%�:�K���&����A��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����c��X
�����4�&�2�u�%�>���T���F��1�����
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�K����Z	��G��U��4�
�:�&��+�E��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�0�<�3�<�(���P����[��=N��U���u�u�u�u�w�}�W���&����\��E��I���
�
�0�<�3�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�0�4�6���������@��YN�����&�u�x�u�w�-�B�������l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�b�?����	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�<�(���&����Q�����ߊu�u�u�u�w�}�W���Y���F��1�����%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W���Y�Ʃ�@�������7�1�c�|�#�8�W���Y���F�N��U���u�u�u�
��8����&����C��R�����7�!�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����7�!�
�'�0�<����Y����V��C�U���%�`�7�!��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h�����0�u�h�4��2�����ԓ�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
��8����&����O��_�����u�u�u�u�w�}�W���Y����Q��h����u�
�
�0�6�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���&�<�;�%�8�8����T�����T��U´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������W������u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$�������^9����U���}�4�
�:�$�����&���T��Q1�����3�
�f�
�'�9����P�Ƹ�VǻN��U���u�u�u�u��3��������e+��G������
�
�
�2��E���DӁ��l ��h��*���d�g�4�
�2�(���s���F�N��U���3�
�:�0�#�/�(���8����q��d)�����'�2�g�e�k�}����&ù��9��h_�*���'�!�'�
�l�}�W���Y���F������
�0�8���1��������l��R	��G���h�2�%�3�g�;�F���&����R��R����_�u�u�u�w�}�W���Y����\��C��*����%�4�0�6��(�������F�	��*���
�
�
� �f�o��������lU��N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y����[��R�����0�}�%���.�^ϱ�Y����@��RN�����0�u�x�u�w�<�(�������@��Y1�����u�'�6�&�w�<�(������R��RB�����2�7�1�l�{�:����I����l ��]�����:�0�u�'���(���&����T��G1�����u�u�7�2�9�}�W���YӅ��VF��h-�����<�_�u�u�w�}�W�������C9��h��*���
�u�k�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���&�2�7�1�n�t�^Ϫ����F�N��U���u�u�u�4������E�ƭ�l5��D�����d�_�u�u�w�}�W���Y�Ʃ�@ǻN��U���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}��������l��h��*���k�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ����F��*���&�
�:�<��}�W���&����U9��Q��F؊�%�1�;�|�~�}����Y���F�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}�W�������F�N��U���u�u�u�u�6��$������R��c1��G���8�d�_�u�w�}�W���Y���V��^�U���u�u�u�u� �8�W���*���� 9��Z1�H���u�u�u�u�w�}�W��������T�����2�6�d�h�6������Ƣ�GN��G1�����9�2�6�e�j�:����I����l ��Z�����:�0�|�|�#�8�}���Y���F�N��U���4�
��3�:�a�W���*����9��Z1����u�u�u�u�w�}�W������F�N��U���u�u�u�%������DӇ��`2��C]�����n�u�u�u�w�}�W���YӃ����=N��U���u�u�u�=�9�2����Y���9F�N��U���u�u�u�%������D�Ĕ�kD��N��U���0�1�6�&�l�}�Wϻ�Ӗ��P��dךU���x�4�
�:�2�<����Y����V��C�U���4�
�:�0�6�.���������T��]���6�y�2�%�1�m��������9��h
�����%�&�2�6�2��#���J����lT�N�����;�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$�������^9����U���}�4�
�:�$�����&���T��Q1�����3�
�a�
�'�9����P�Ƹ�V�N��U���u�u�4�
�8�8�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���%�<�9�u�$�4�Ϯ�����F�=N��U���<�9�
�&�>�3����Y�Ƽ�\��DF��*���'�y�4�
�>�����*����9��Z1����u�0�<�_�w�}�W�������\�V�����
�:�<�
�w�}���������F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�|�#�8�W���Y���F������u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����VF������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��R��U���<�;�%�:�2�.�W��Y����C9��V
�����2�
�'�6�m�-����
ۇ��P�P�����3�g�3�
�c���������C9��P1������&�f�3�:�o�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ�ӈ��N��h�����:�<�
�u�w�/�(���&����U��\�����;�|�|�u�?�3�}���Y���F�V�����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����W�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����D�����d�e�4�&�0�}����
���l�N��*���
�1�
�d��.����	����	F��X��´�
��3�8�]�}�W������F�N��U���u�4�
�<��9�(��Y���R��X ��*���
�u�u�%������Y����G	�G�U���0�1�%�:�2�.�}�ԜY�����D�����d�d�4�&�0�}����
���l�N��*���
�1�
�c��.����	����	F��X��´�
��3�8�]�}�W������F�N��U���u�4�
�<��9�(��Y���R��X ��*���
�u�u�%������Y����G	�G�U���0�1�%�:�2�.�}�ԜY�����D�����d�d�4�&�0�}����
���l�N��*���
�1�
�b��.����	����	F��X��²�%�3�e�3�e�;�(��&����\�������6�0�
��$�n����K���F��P��U���u�u�u�u�w�}��������W9��N�U���%�6�;�!�;�:���DӇ��@��T��*���&�f�3�8�e�}��������C9��Y�����6�e�h�2�'�;�G���K����R��V�����|�n�u�u�2�9��������9l�N�U���&�2�7�1�f�}����Ӗ��P��N����u�%�&�2�5�9�Fց�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������Z���6���&�}�u�:�9�2�G���Y����\��h��*���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�b�6�.��������@H�d��Uʴ�
�<�
�1��j��������\������}�%�&�4�#�}��������B9��h��*���
�y�%�e�6�-����&����9F����ߊu�u�u�u�w�}�W���	����l��h]�I���}�%�6�;�#�1����H����lV��[��*���#�1�u�;�w�2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��\�ߊu�u�;�u�%�>���s���K�V�����1�
�c�4�$�:�W�������K��N�����<�
�1�
�a�<����&����\��E�����%�&�4�!�w�-��������`2��C_�����y�%�d�8�/�<�(���P�����^ ךU���u�u�u�u�w�}��������lR��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�l��������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*���4�&�2�u�%�>���T���F��h��*���
�`�4�&�0�����CӖ��P�������!�u�%�&�0�>����-����l ��h^�����'�:�
�'�+��ԜY�Ʈ�T��N��U���u�u�u�u�6���������Z� ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
��8��������WO�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��4�&�2�u�%�>���T���F��h��*���
�m�4�&�0�����CӖ��P�������!�u�%�&�0�>����-����l ��h^����7�!�
�%�!�9�}���Y����]l�N��U���u�u�u�4��4�(���&���F��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
�2�<�������9F���U���6�&�n�_�w�}�Z���	����l��hW����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*���4�&�2�
�%�>�MϮ�������D�����
�
�9�=��-��������TJ��h_�����%�#�1�<��4�[Ϯ�K����Z	��V�����;�&�2�u����������W9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�l�u�h��-�B�������l��h�����h�4�
�:�$�����&����AF��h\�����1�4�
�9��3����DӇ��P	��C1�����e�u�'�}������	����l��D��Hʴ�
�:�&�
�8�4�(�������lV��[��*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�4�
�!�%�}�W�������l
��^��\��u�u�0�1�'�2����s���F������6�0�
��$�l����IӇ��Z��G�����u�x�u�u�6�����
����g9��1�����4�&�2�
�%�>�MϮ�������D�����d�|�u�u�5�:����Y����������7�1�d�|�#�8�W���Y���F������6�0�
��$�l����I���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�&�2�6�2��#���H����lV�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����D�����
��&�g�1�0�FϿ�
����C��R��U���u�u�4�
�>�����*����9��Z1�����2�
�'�6�m�-����
ۇ��@��U
��D��_�u�u�0�>�W�W���Y�ƥ�N��h��*���
�d�|�!�2�}�W���Y���F��G1�����0�
��&�e�;���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�f�3�:�o�����Ƽ�\��D@��X���u�4�
�<��.����&����U��1�����
�'�6�o�'�2��������T9��S1�D�ߊu�u�0�<�]�}�W���Y���R��^	�����c�|�!�0�w�}�W���Y�����D�����
��&�f�1�0�E��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�D������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӁ��l ��h��*���d�g�4�
�2�<����Y����V��C�U���2�%�3�e�1�l����J����l��V�����'�6�o�%�8�8�ǿ�&����P��h=�����3�8�e�u�'�>�[Ͽ�&����Q��\����<�
�&�$���݁�
����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u�_�������l
��^��U���%�&�2�6�2��#���H����lV�V �����4�
�<�
�3��E�������C9��Y�����6�d�h�4��4�(�������@��Q��D���|�!�0�u�w�}�W���Y����A��h^��*ۊ� �d�g�4��8�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F�	��*���
�
�
� �f�o�������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}�����֓�lW��B1�G���
�!�'�u�j�:����I����l ��]�����!�'�
�%�$�<�������F��G1��E���d�3�
�f��3�������F��1�����<�
�<�n�w�}�����֓�lW��B1�G���
�0�4�e�k�}�(ځ�����]9��PUךU���'�
�
�
�����K����^��N�U���
�4�
�;�$�:�}���Y���T��Q1�����3�
�a�
�'�>�W�������A	��D�X�ߊu�u�'�
���(݁�����l��T�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�e�;���Y����U9��Q1�����f�
�%�1�9�q��������V��c1��F���8�g�_�u�w�8��ԜY���F��F�����:�&�
�:�>��W���	������F�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9����Q����\��h�����u�u�'�
���(ށ�����l��S��\���:�u�4�
�8�.�(�������F��h��*���$��
�!��.�(���P�Ƹ�V�N��U���u�u�2�%�1�m��������9��h��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�:����I����l ��Z�����0�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]ǑN�����3�e�3�g�1��C݁�	����A�
N�����e�3�g�3��i�(���
����l��D�����2�_�u�u�%��(߁�&����lW��h��%���:�
�u�h�'�o�'�������l��d��Uʲ�%�3�e�3�e�;�(��&����C��R ��E��u��;�1��8����4����R$��V=��*���0�
�g�n�w�}�����֓�lT��B1�G���
�%�'�0�#�l�K���*����V9��E��#���%�4�0�4���(ށ�����]ǻN�����
�
�
�
�"�l�E���&����P��h\��Hʳ�
�:�0�!�%��!���	����G��{1��G���2�g�e�_�w�}�Z���&ù��C��V�����;�&�2�4�$�:�W�������K��N�����4�%�4�4��1�(���
����@��Y1�����u�'�6�&���(�������l��N��E���%�4�4�
�;�����s���Q��Yd��U���u�<�u�}�'�>��������lW���*���=�
�%�#�3�t����Y���F�N��U���
�9�=�
�'�+����&����[��h^�����
�%�#�1�]�}�W���Y����l�N��U���u�%�e�4�'�<��������l��R�����4�%�4�4��1�(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����4�%�4�<��4�W�������A	��D�X�ߊu�u�
�
�;�5�(���
����@��Y1�����u�'�6�&���(�������lV��[��*���2�u�
�
�;�5�(������F�U�����u�u�u�<�w�u��������\��h_��U���
�9�=�
�'�+��������9F�N��U���u�
�
�9�?��������C9��V���ߊu�u�u�u�;�8�}���Y���F�G1�����4�<�
�<�w�`��������l��PUךU���u�u�;�u�1�}�W�������A	��D����u�
�`��4�2�W������W��R��&���9�=��!����������lǻN��Xʥ�d�
�0�!�%�<�(���Y����T��E�����x�_�u�u��h�$�������l��h�����%�:�u�u�%�>����	������h��*���
� �d�g�6�����Y����Z��D��&���!�
�&�
�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�f�3�8�e�}��������C9��Y�����6�e�h�2�'�;�G���K����R��V�����|�|�!�0�w�}�W���Y�����1�����
�%�#�1�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����1�����
�%�#�1�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�f�0����&����Z��^	�����;�%�:�0�$�}�Z���YӖ��l��h�����<�
�<�
�$�4��������C��R�����8�-�4�
�;�q��������C9��S1�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���&����_����ߊu�u�u�u�w�}�(ށ�����l��h�����i�u�
�
�6��������F�N�����u�u�u�u�w�}��������C9��S1��*���u�h�%�d�:�%��������V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�%�d�8�/�4�(���Y����T��E�����x�_�u�u����������l��^	�����u�u�'�6�$�u�(ށ�����lW��V�����u�
�
�4��-����s���Q��Yd��U���u�<�u�}�'�>��������lW���*���
�%�#�1�~�)����Y���F�N��*ۊ�4�
�;�&�0�a�W���&����9F�N��U���0�_�u�u�w�}�W���&¹��K9��h��U��%�d�8�-�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��h\�����1�4�
�9��3��������]F��X�����x�u�u�%�e�����&����_��Y1�����&�2�
�'�4�g��������lT��R�����
�9�y�%�e�����&����_��E�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�e�����&����_����ߊu�u�u�u�w�}�(݁�����l��A�����<�u�h�%�e�����&����_��N��U���0�&�u�u�w�}�W���YӖ��l6��^�����9�
�;�&�0�a�W���&����\��G1�����0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�K����Z	��^ �����&�<�;�%�8�8����T�����h>�����<�
�<�
�$�4��������C��R������'�:�y�'�o�'�������V�G1��%���:�
�%�#�3�W�W�������F�N�����}�%�6�;�#�1����H����lT��R�����
�9�|�u�?�3�}���Y���F�G1��%���:�
�;�&�0�a�W���&����\��N��U���0�&�u�u�w�}�W���YӖ��l6��^�����<�u�h�%�e�����&����l�N��Uʰ�1�<�n�_�w�}��������@]ǑN����� ��8�;���W������lV��h\�� ��g�4�
�0�"�3�G�ԶY���F��1��!���;�
�
�
�'�+�Ͽ�
����C��R��U���u�u�%�a��	����&����R��[
�����;�%�:�u�w�/����Q����VJ��E��*ڊ�
�
� �d�e�<�(����ƭ�l��h�����
�!�
�&��t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�f�3�:�o�W���Y������T�����2�6�e�h�0�-�����ԓ�F9��1��*���0�|�|�!�2�}�W���Y���F��hZ��*���<�2�0�e�6�����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N����� ��8�;���(������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�}�WϮ�M����Z��P1��D��u�'�
�
���(���H�ԓ�C9��C��*��_�u�u�x�'�i�"�������V9��V�����&�<�;�%�8�8����T�����h;�����2�0�d�4��1�(�������A	��N�����&�4�
�0�w�/�(���&����U��\�����;�y�4�
�>�����*���� 9��Z1����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GU��D��\ʴ�1�;�!�}�'�>��������lV�	��*���
�
�
� �f�o�������O��_�����u�u�u�u�w��(�������l��h�����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϮ�M����Z��P1��D���
�9�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�2�<��������l�������%�:�0�&�w�p�W���	�ӓ�V��V�����;�&�2�4�$�:�(�������A	��D��*ߊ�0�4�4�
�;�q��������R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�B�������l��G�����_�u�u�u�w�}�W���&����l��A�����<�u�h�%�b�?����	����l�N��Uʰ�&�u�u�u�w�}�W���	�ӓ�V��V�����;�&�2�i�w��(�������E
��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�h����&����Z��D��ʥ�:�0�&�u�z�}�WϮ�L����R9��h��*���<�;�%�:�w�}����
�μ�9��C����7�!�
�'�0�}�(ځ�����C9��SGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�`�5�)�(��������YNךU���u�u�u�u����������TF���*���4�_�u�u�w�}����s���F�N�����7�!�
�;�$�:�K���&ƹ��G��E�����u�u�u�;�w�;�W���YӃ����T��N�ߊu�u�
�
��4�������F��G1��E���g�3�
�a��-��������9l�N�U���
�
�<�<�0�8�G���&����R��P �����&�{�x�_�w�}�(ف�&����]��h^�����1�4�&�2��/���	����@��G1��Yʲ�%�3�e�3�e�;�(��&����\�������6�0�
��$�n����K���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�(���&����]��X�����:�&�
�:�>��W�������9��1��*��
�%�1�;�~�t�W������F�N��Uʥ�c���8�9��(߁�	����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�
�
��4�����֓�C9��SN�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���C9��a1�����
�
�u�h�0�-�����ԓ�F9��1��*��� �;�f�_�w�}�Z���&Ź��g��Y	��*ۊ�%�#�1�4�$�:�W�������K��N�������8�;���(�������@��Y1�����u�'�6�&��-�������lV��h\�� ��g�4�
�:�2�}��������B9��h��*���
�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��F���8�g�u�;�w�2�_ǿ�&����G9��P��E��2�%�3�e�1�o����M����l��RG��\ʡ�0�u�u�u�w�}�W���	�Г�l2��^ �����4�
�9�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���C9��a1�����
�
�
�%�!�9�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�u�u�%�o�
��������F�	��*���
�
�
� �f�o��������lR��=N��U���%�m��!�:�3�(���&����_��D��ʥ�:�0�&�u�z�}�WϮ�A����Z��P1��E���
�9�
�&�>�3����Y�Ƽ�\��DF��*���u�'�
�
���(���H�ԓ�C9��Y����<�
�&�$���܁�
����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������F��SN�����%�6�;�!�;�:���DӁ��l ��h��*���d�g�4�
�8�8�^�������9F�N��U���u�
�
�
�>�4����I����E
��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�%�o�
��������9��h��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƹF��hV��*���<�2�0�d�k�}����&ù��9��h_�*���'�!�'�
�l�W�W���TӖ��l1��^�����d�4�
�9�w�.����	����@�CךU���
�
�
�<�>�:��������W9��D��*���6�o�%�:�2�.�����ƫ�C9��1��G���
�a�
�%�3�3�[Ͽ�&����P��h=�����3�8�g�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9����Q����\��h�����u�u�'�
���(݁�����l��S��\���u�=�;�_�w�}�W���Y�Ƽ�9��C�����
�
�%�#�3�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��hV��*���<�2�0�d�6�����DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�;�w�8���