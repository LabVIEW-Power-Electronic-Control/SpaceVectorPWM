-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ��m�d�a��}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e�4�%�4�m��W���&����p9��t:��U��u�:�;�:�g�f�W�������\��yN��1�����_�u�w��(�������l��T��;ʆ�����]�}�W���&����	F��=��*����
����u�FϺ�����O��N�����8�-�4�
�;�}�W���*����|!��d��Uʥ�g��'�:�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����c��X
�����1�o��u���8���B�����h;�����2�0�e�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���&ǹ��g��Y	��*ڊ�%�#�1�o��	�$���5����l�N��A����8�;�
��}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y����lR��h:�����0�d�4�
�;�}�W���Y����)��tUךU���
�
�0�4�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ӓ�V��V�����u������4�ԜY�Ƽ�9��c�����
�u�u� �w�	�(���0����p2��F�U���;�:�e�n�w�}����/����Z��R1�����9�u�u� �w�	�(���0��ƹF��hX��*���<�2�0�d�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����e9��Z��*���
�%�#�1�m��#ύ�=����z%��N������!�8�;���W���,�Ɵ�w9��p'��#����u�f�u�8�3���B�����h9�����2�0�e�4��1�W���,�Ɵ�w9��p'�����u�
�
�
�>�4����H����f2��c*��:���
�����l��������l�N��M���!�8�;�
����������f2��c*��:���u�n�0�1�]�W��������A��R��U���8��m�d�c��W���s���R��^��ʖ��
�����9���?����`2��y)�U���4�!�<� �2��%���<����g/��h'��:ʺ�u�0�4�u�w�/����������N��W���m�d��3�g�5����&����lR��"��<������h�/�q�;���7����u*��cS�=���������GÖ�*����f2��v<�����e�e�9�a�c�l�?���0����l%��t%��@��e�e�y����"���+����G��DB��&�������e�s�O��I߮��l5��h"��H�������	����U����`?��z+��EƝ������l�[���&����u �\�=�������o�n�
��Y����\��V �����:�&�
�:�>��W���-����t/��S��D��u�u�6�;�#�3�W�������l
��^��U����
���w�`�P���s���P	��C��U����
�!�
�$��W���-����t/��a+��:���g�1�"�!�w�t�M���I���9F������!�4�
��$�o����H����g"��x)��*�����}�u�8�3���Y���W��d��Uʶ�;�!�;�u�'��(���&����F��d:��9�������w�o��������\�_�W�ߊu�u�:�&�6�)��������_��h^��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�:�$�<�Ͽ�&����G9��1�Oʆ�������8���Iӂ��]��G��H���w�_�u�u�8�.��������]��[�*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�d�w�_�w�}�����ƭ�l%��Q��Oʆ�������8���Kӂ��]��G��H���e�w�_�u�w�)�����ƪ�^9��T�����u�!�<�2�]�}�W�������VF��Z1�����;�u�3�4������Cӕ��]��^�����w�_�u�u�>�3�Ͽ�&����P��h=�����3�8�e�o���;���:���F��P ��U���&�2�7�1�f�}�W���5����9F������%�e�4�%�6�4�(���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����4�%�4�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���@��V��*ڊ�9�=�
�%�!�9��������`2��{!��6�ߊu�u�<�;�;�-�G���	����C9��S1�����u��
���}�J���^���F��P ��U���
�4�
�;�$�:�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��h_�����'�2�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�e�l�}�Wϭ�����C9��Z�����9�
�;�&�0�g�$���5����l�N�����u�
�
�4��-����	����	F��s1��2���o�u�e�n�w�}�����Ƽ�9��E��*���&�2�o����0���/����aF�N�����u�|�_�u�w�4����	�ԓ�V��S1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�ԓ�V��S1��*���
�;�&�2�m��3���>����F�D�����
�
�0�<�3�<�(���&����\��c*��:���u�h�r�r�]�}�W�������lS��R�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&ƹ��G��E��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��n�u�u�&�0�<�W���&����l��A�����<�u�u����>��Y����Z��[N��@���!�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���
����W��N�7�����_�u�w�4��������W��R��&���9�=��!����������\��c*��:���
�����l��������l�N�����u�%�&�2�4�8�(���
�ԓ�@��T��!�����n�u�w�.����Y����Z��S
��E���u����l�}�Wϭ�����T��Q1�����3�
�g�
�'�9����Y����)��tUךU���<�;�9�3��2��������~'��_������&�d�'�0�o�G��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������
�0�8���1��������l��h��*��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����U9��Q��Gۊ�%�&�4�!�m��3���>����F�D�����'�
�
�
�����H����Z��T��!�����n�u�w�.����Y����U9��Q1�����g�
�%�'�6�$�Mύ�=����z%��N�����4�u�'�
���(ށ�����l��V����o������!���6���F��@ ��U���_�u�u�<�9�1�����֓�lW��B1�D���
�4�
�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��1��D���
�g�
�;�5�)�(���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����e�3�d�3��o�(�������]9��N��1��������}�D�������V�=N��U���;�9�2�%�1�m��������9��h�� ���d�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����l ��h��D���4�
�0� �9�o�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E��*ڊ�
�
� �d�f�<�(���Cӵ��l*��~-�U���&�2�4�u�%��(߁�&����lW��h�����!�o�����4�ԜY�ƿ�T��	��*���
�
�
� �f�l�������5��h"��<��u�u�&�2�6�}����&ù��9��h_�*���<�9�u�u���8���B�����Y�����3�e�3�g�1��Dށ�	����W�=��*����n�u�u�$�:��������9��1��*��
�;� �0�4�3�(���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����e�3�g�3��n�(���)����W9��N��1��������}�D�������V�=N��U���;�9�2�%�1�m��������9��h8�����!�d�o����0���/����aF�N�����u�|�_�u�w�4��������lV��h\�� ��d�<�
�%�%�8���Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
�
�
�
�"�l�F���&����A��T��!�����
����_������\F��d��Uʦ�2�4�u�'���(���&���� W��G1�����
�u�u����>���<����N��
�����e�n�u�u�$�:��������9��1��*��
�%�'�!�%��W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����3�g�3�
�d��������� F��d:��9�������w�n�W������]ǻN�����9�2�%�3�g�;�E���&����R��R����o������!���6���F��@ ��U���_�u�u�<�9�1�����֓�lT��B1�D���
�0� �;�b�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��*���
� �d�d�6����*����|!��d��Uʦ�2�4�u�%�$�:����&����GU��D��U����
���l�}�Wϭ�����R��^	�����`�u�u����L���Yӕ��]��P�����3�d�3�
�e���������C9��V�����o������M���I��ƹF��^	��ʲ�%�3�e�3�e�;�(��&����G��h�����!�'�2�o���;���:���V�=N��U���;�9�4�
��;���*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V�����1�
�b�o���2���s���@��V�����2�7�1�d�`�g�5���<����F�D�����%�&�2�7�3�i�W���6����}]ǻN�����9�4�
�<��9�(��CӤ��#��d��Uʦ�2�4�u�%�$�:����O����q)��r/�����u�6�8�:�2�)�ݚ�A�׈�U9��Q1�<�ߊu�u�:�!��}�W���YӇ��P
��N��U���
���n�w�}�W�������GF��~ ��!�����n�u�w�}�WϿ�&����GF��~ ��!�����n�u�w�}�WϿ�&����\��b:��!�����n�u�w�}�WϿ�&����\��b:��!�����n�u�w�}�WϿ�&����JF��x;��&������_�w�}�W�������[��T��;ʆ�������8���J�ƨ�D��^����u�u�u�;�:�%�E��0�Ɵ�w9��p'��#����u�f�u�8�3���B���F������
�u�u����;���:����g)��]����!�u�|�_�w�}�W���	����F��N�:���������4���Y����W	��C��\�ߊu�u�u�u�'�/����&����|3��d:��9�������w�n�W������]ǻN��U���%�'�!�'��}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y���F��G1��U���������^�ԜY�Ʃ�WF��Z�����_�_�u�u�8�-����Y�Ԉ�W����*���u��u�u�'�/�W�ԜY���F��h��U���������}���Y���R��D��U��������W�W���Y�ƭ�l��E��U��������W�W���Y�ƭ�l��RN�:��������W�W���Y�ƭ�l��RN�:��������W�W���Y�ƭ�l��S��U���u��
���f�W���Y����]9��R�����u�u�����0���/����aF�N�����u�|�_�u�w�}�W���)����W9��N��U���
���
��	�%���Hӂ��]��G�U���u�u�<�
�'�/����H����}F��s1��2������u�d�}�������9F�N��U����0�6�;��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY���F��h�� ���e�o�����;���:����g)��]����!�u�|�_�w�}�W���	����F��N�:���������4���Y����W	��C��\�ߊu�u�u�u�'�/����&����|3��d:��9�������w�n�W������]ǻN��U���%�'�!�'��}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y���F��G1�����
�u�u� �w�	�(���0����p2��F�U���;�:�e�n�w�}�W�������G��h[��U���u��
����2���+������Y��E��u�u�u�u�6����0�Ɵ�w9��p'��\�ߊu�u�;�u�8�-����B��ƓQ��Yd��Uʲ�%�3�e�3�f�;�(��Y�Ư�^��R ��ؑ�m�d�a�
���}���Y������FךU���u�u�%�6�<�`�W�������F�N�����&�u�k�4��.�[���Y�����D����u�'�
�
���(���H�ד�C9��V�����u�u�u�%�3�3�W�������lV��h_�� ��d�4�
�:�2�W�W���Y�ƭ�l��RN��U���
�
�
�
��(�F�������_�N��U���4�
�0�1�w�c�����֓�lW��B1�D���
�0�1�y�w�}�W�������C��N��U���
�
�
�
��(�F�������C��BךU���u�u�;�8�/�o�J�������9��1��*��
�;�8�-�e�W�W���Y�ƥ�l��V1�H���'�
�
�
�����H����Q��h^�U���u�u�4�
�2�(���D�ƫ�C9��1��D���
�g�
�%�%�)����U���F������'�
�u�k�0�-�����ד�F9��1��*��� �;�d�_�w�}�W���	����F��N��U���
�
�
�
��(�F�������G��h\�U���u�u�4�
�2�`�W���&����U9��Q��Gۊ�%�6�|�_�w�}�����֓�lT��B1�D��6�8�:�0�#�0�3��H�Ҫ�9��d��Uʥ�'�u�4�u�]�}�W���Y����_�	N��*���y�u�u�u�w�<�(���Y����C9��CBךU���u�u�%�&�6�)�J�������9��1��*��
�%�&�4�#�W�W���Y�ƭ�l��RN��U���
�
�
�
��(�F�������]�N��U���4�
�1�0�j�}����&ù��9��h_�*���<�9�y�u�w�}�WϿ�&����JF�	��*���
�
�
� �f�l��������9F�N��U��� �0�6�;��}�IϹ�	����l ��h��D���<�
�%�'�2�)�G�ԜY���F��h>�����f�h�u�'���(���&���� W��Y1�����
�y�u�u�w�}����	����]��S����3�e�3�g�1��Dށ�����A��C1����u�u�u�;� �8����&�����h��*���
� �d�d�>���������l�N��Uʴ�
�0� �;�g�`�W���&����U9��Q��Fۊ�%�'�!�'��q�W���Y����C9��C��*���k�2�%�3�g�;�E���&����R��R����_�u�u�u�w�-��������X��E��*ڊ�
�
� �d�f�<�(�������l�N��Uʴ�
�0� �;�d�`�W���&����U9��Q��Fۊ�%�'�!�'��q�W���Y����C9��C��*���k�2�%�3�g�;�E���&����R��R����_�u�u�u�w�-��������X��E��*ڊ�
�
� �d�f�<�(�������l�N��Uʴ�
�0�h�u�%��(߁�&����lW��h�����_�_�_�u�w�p�W���Y����V��D�����%��
�&�~�2�W���Y����VF��T�����x�u�u�4����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��G1��*���u�h�4�
��.�F�������F�N��U���0�&�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��=N��U���u�u�u�u�w�}�W���:����^F���;���&�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�P�����3�d�3�
�e���������C9��V�����4�&�2�u�%�>���T���F��G1��E���d�3�
�g��-��������@��C1�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�2�'�;�G���H����T��V�����
�%�&�4�#�/���Y����\��h�����n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}����PӇ���������7�1�l�|�~�)����Y���F�N��U���u�u�'�
���(ށ�����l��D�����
�!�'�
�2�}�JϿ�&����G9��P��D�ߊu�u�u�u�w�}�W�������N��h�����:�<�
�u�w�/�(���&����U��_�����4�,�|�!�2�}�W���Y���F�N��U���'�
�
�
�����H����@��C1��*���'�
�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W������lV��h\�� ��d�4�
�!�%���������V��D��ʥ�:�0�&�u�z�}�WϹ�	����l ��h��D���4�
�!�'��-��������l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�
�
�
��(�F�������R��V�����
�0�u�h�6�����&����P9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���g�3�8�d�w�3�W���Qۇ��P	��C1�����e�h�2�%�1�m��������9��h
�����|�!�0�u�w�}�W���Y���F�N�����
�
�
�
�"�l�F���&����G9��h�����0�u�h�4��2��������]ǻN��U���u�u�u�u�;�4�W���	����@��X	��*���u�'�
�
���(���H�ד�C9��V
��\ʡ�0�u�u�u�w�}�W���Y���F��E��*ڊ�
�
� �d�f�<�(�������l��E�����h�4�
�:�$�����&��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m��������E
��G��U���<�;�%�:�2�.�W��Y����lV��[��*���#�1�%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����R
��V1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�0�$�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���Yӏ����D�����d�b�u�=�9�W�W���Y���F�N��U���u�%�e�4�'�<��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&���G��d��U���u�u�u�u�w�}�W���YӖ��l��_�����1�%�0�u�j�-�G���	����C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(߁�����C�������%�:�0�&�w�p�W���	�֓�_��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�g�<����	����[��G1�����9�f�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʥ�e�4�%�4�6���������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�~�)����Y���F�N��U���u�u�
�
�;�5�(������C9��V���ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lW��V�����1�%�0�u�$�4�Ϯ�����F�=N��U���
�4�
�%�!�9����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����2�7�1�d�`�}����s���F�N��U���u�u�u�u�'�l��������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&����P�C��U���u�u�u�u�w�}�W���Y�����h��*���#�1�%�0�w�`��������C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(ށ�����V��D��ʥ�:�0�&�u�z�}�WϮ�H����l��P1�����
�'�6�o�'�2��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�u�f�t����s���F�N�����4�
�&�u�w�l�^Ϫ����F�N��U���u�%�d�8�/�-����DӇ��P	��C1��F؊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����^��V�����|�!�0�u�w�}�W���Y���F�N��*ۊ�4�
�'�2�k�}�(ށ���ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�o�'�������l��h��ʴ�&�2�u�'�4�.�Y��s���C9��g�����%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��E��*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z �V�����1�
�c�|�#�8�W���Y���F�N��U���u�u�u�
��8��������W9��R	��Hʴ�
�:�&�
�8�4�(��Y���F�N��U���u�u�9�<�w�<�(���&����S�C��U���u�u�u�u�w�}�W���Y�����h>�����4�
�9�
�%�:�K���&����A��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����c��X
�����4�&�2�u�%�>���T���F��1�����
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�K����Z	��G��U��4�
�:�&��+�E��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-��������\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�0�<�3�<�(���P����[��=N��U���u�u�u�u�w�}�W���&����\��E��I���
�
�0�<�3�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�0�4�6���������@��YN�����&�u�x�u�w�-�B�������l��h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�b�?����	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�<�(���&����P�����ߊu�u�u�u�w�}�W���Y���F��1�����%�#�1�%�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W���Y�Ʃ�@�������7�1�c�|�#�8�W���Y���F�N��U���u�u�u�
��8����&����C��R�����7�!�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����7�!�
�'�0�<����Y����V��C�U���%�`�7�!��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h�����0�u�h�4��2�����ԓ�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
��8����&����O��_�����u�u�u�u�w�}�W���Y����Q��h����u�
�
�0�6�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���&�<�;�%�8�8����T�����T��U´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������W������u�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$�������^9����U���}�4�
�:�$�����&���T��Q1�����3�
�g�
�'�9����P�Ƹ�VǻN��U���u�u�u�u��3��������e+��G������
�
�
�2��F���DӁ��l ��h��*���d�d�4�
�2�(���s���F�N��U���3�
�:�0�#�/�(���8����q��d)�����'�2�g�`�k�}����&ù��9��h_�*���'�!�'�
�l�}�W���Y���F������
�0�8���1��������l��R	��E���h�2�%�3�g�;�F���&����R��R����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9F�C����;�-�u�!�#�}����*����F����U���!�u�4�=�9�s�Z�ԜY�ƭ�l(��Q�����2�
�'�6�m�-����
�έ�l%��Q��U���6�y�4�
�>�����I�ƫ�C9��1��D���
�g�
�%�3�3�[Ϲ�	����l ��h��D���4�
�:�0�]�}�W������F�N�����%��
�&�w�.�W���Y���F��_������&�d�3�:�m�J���Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�;�!�4��4�(���&���F��R ךU���u�u�u�u�w�}�W���	����U��S�����
�!�
�&��f�W���Y���F�N�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�f�;���s���F�N��U���0�1�<�n�w�}�W���Y����[��V��!���g�3�8�d�j�}�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�}�%�6�9�)���������h��*���
� �d�d�6�����P����[��N��U���u�u�u�u�w�}����*����Z�V��!���f�3�8�g�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:��ي�&�
�u�k�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����4�
�:�&��2����Y�ƫ�C9��1��G���
�f�
�%�3�3�^���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:��ۊ�&�
�n�u�w�}�W���Y�����Rd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�f�3�8�e�W�W���Y���F�N��ʼ�n�u�u�u�w�}�Wϩ��ƣ�[��S�U���u�u�u�u�w�}�WϿ�&����@�
N��-���_�u�u�u�w�3�W������F��SN�����&�_�u�u�z�}�����ƭ�@�������{�x�_�u�w�-����&����T��E��Oʥ�:�0�&�4��8�W���&����U9��Q��Fۊ�%�1�;�y�6�����
����g9��1����_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C]�����|�4�1�;�#�u��������\��h^��U���
�
�
�
��(�F�������]�G�����_�u�u�u�w�}�W�������[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�:�2�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������]F��X�����x�u�u�4��9����
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�|�u�w�?����Y���F��QN�����}�%�6�;�#�1����H����C9��V��\ʴ�1�}�%�6�9�)���������D�����
��&�d�1�0�G���Y����l�N��U���u�4�
�1�2�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���'�4�,�4�$�:�W�������K��N�����0�1�
�&�>�3����Y�Ƽ�\��DF��*���u�'�
�
���(���H�ד�C9��Y����<�
�&�$���܁�
����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������F��SN�����%�6�;�!�;�:���DӁ��l ��h��*���d�d�4�
�8�8�^�������9F�N��U���u�%�'�4�.�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��m�W�������A	��D�X�ߊu�u�%�&�0�?���A����Z��G��U���'�6�&�}�'��(���P�����^ ךU���u�u�u�u�w�}��������lW��R��]���6�;�!�9�f�l�JϿ�&����@�
�����d�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��h�W�������A	��D�X�ߊu�u�%�&�0�?���O����Z��G��U���'�6�&�}�'��(���P�����^ ךU���u�u�u�u�w�}��������lW��R��]���6�;�!�9�f�l�JϿ�&����@�
�����g�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��k�W�������A	��D�X�ߊu�u�%�&�0�?���N����Z��G��U���'�6�&�}�%��(߁�&����lW��h�����y�4�
�<��.����&����U��GךU���0�<�_�u�w�}�W���Y���R��^	�����c�u�h�}�6�����&����P9��
N��*���
�&�$���)�(���&����]��X�����:�&�
�:�>��W�������9��1��*��
�%�1�;�~�t�}���Y����C��R���ߊu�u�x�4��4�(���&����@��YN�����&�u�x�u�w�<�(���&����_��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��L��u�4�
��1�0�GϺ�����O������!�9�d�d�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���Y����T��E�����x�_�u�u�'�.��������R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���&����R9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�f�u�h��<�(���
����T��N�����4�%�4�4��1�^Ͽ�ӈ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�6�����&����P9��
N��*���'�|�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�C���
������T��[���_�u�u�%�$�:����MŹ��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(ށ�����l��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����^��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�`�w�.����	����@�CךU���%�&�2�7�3�h�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�u�
��8��������WOǻN�����_�u�u�u�w�}�W���Y����Z��S
��@��u�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�K����Z	��V�����n�u�u�0�3�-����
��ƓF�C�����2�7�1�c�w�.����	����@�CךU���%�&�2�7�3�k�(�������A	��N�����&�4�
�!�%�q��������V��c1��D���8�e�u�
��8����&����9F����ߊu�u�u�u�w�}�W���	����l��hX�I���;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`��������R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�l�u�&�>�3�������KǻN�����2�7�1�l��.����	����	F��X��´�
�!�'�y�'�m��������E
��^ �����%�d�8�-�6���������F��1�����
�%�#�1�>����	�ӓ�V��V�����;�&�2�_�w�}����s���F�N��U���4�
�<�
�3��G��Y�μ�9��C�����1�<�
�<�w�}��������\��h^�����%�g��'�8���������@��
N��*���&�
�:�<��t����	�ד�R��G1�����
�<�u�u�'�>��������lV�X�����4�%�4�4��1�(���
�����T�����2�6�e�u�%�u���������T�����2�6�e�|�]�}�W���Y����V��=dךU���x�4�
�<��.����&����U��N�����u�'�6�&�y�p�}���Y����Z��D��&���!�
�&�
��.����	����	F��X��´�
�<�
�1��d�}���Y����]l�N��Uʼ�u�4�
�<��9�(��Y����l�N��U���u�4�
�<��.����&����U��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����
����g9��1����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�&�&��(���&����F��D��U���6�&�{�x�]�}�W���
����@��d:��؊�&�
�
�&�>�3����Y�Ƽ�\��DF��*���
�1�
�e�~�}�Wϼ���ƹF�N�����%�&�2�7�3�l�O������F�N��U���4�
�<�
�$�,�$�������^9��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��Q��D��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���܁�
����R��P �����&�{�x�_�w�}��������B9��h��*���
�
�&�<�9�-����Y����V��V�����1�
�`�|�w�}�������F���]���&�2�7�1�f�k�W������F�N��Uʴ�
�<�
�&�&��(���&����F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�4�
�>�����*���� 9��Z1�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N�����e�3�d�3��o�(����ƭ�@�������{�x�_�u�w�/�(���&����U��_�����
�&�<�;�'�2�W�������@N��h��*���$��
�!��.�(������F��h��*���
�e�u�%�$�:����&����GT��D��\���u�7�2�;�w�}�W��������T�����2�6�d�h�6����������T�����2�6�d�h�6�����
����g9��1����u�;�u�:��-��������O�X�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�~�}����s���F�N�����3�e�3�d�1��Eށ�	����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�2�%�3�g�;�F���&����R��RN�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���T��Q1�����3�
�g�
�'�.����E�ƫ�C9��1��D���
�g�
�%�$�<����&����G9��PUךU���'�
�
�
�����H����R
��V1�I���
�
�9�=��3����s���T��Q1�����3�
�g�
�9�?����Y����lS��R�����<�n�u�u�0�-�����ד�F9��1��*���
�u�h�%�f�0����&����9l�N�U���
�
�
�
��(�F���������^	�����0�&�u�x�w�}�����֓�lT��B1�D���
�0�4�&�0�����CӖ��P�������4�
�<�
�$�,�$�������^9��	��*���
�
�
� �f�l�������R��^	������
�!�
�$��^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�}�%�4�3��������[��G1�����0�
��&�e�;���Y����]	�������!�9�2�6�g�`�����֓�lW��B1�D���
�:�0�|�w�/�_�������l
��^��U���%�&�2�6�2��#���J����lT�G�����_�u�u�u�w�}�W���&����U9��Q��Fۊ�%�6�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƫ�C9��1��G���
�f�
�%�4�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�'���(���&���� W��G1�����i�u�'�
���(݁�����l��D�����
�!�'�
�2�f�W�������lV��h\�� ��d�<�
�0�>�9�D��Y����c��X
�����2�_�u�u�%��(߁�&����lW��h�� ���6�;�
�u�j�;�(�������^9��z/�����!���&�%�:�E��s���T��Q1�����3�
�f�
�9���������[��d1�����0�8���;�5�5���*����lW��R	��D��u�u�2�%�1�m��������9��h9�����!�g�i�u��3��������e+��G������
�
�
�2��F��s���K��h^�����
�%�#�1�>�����
������T��[���_�u�u�
��1����	����l��D�����2�
�'�6�m�-����
ۖ��l��_�����1�u�
�
�;�5�(�������A��=N��U���<�_�u�u�w�}��������]��[����h�%�e�4�'�<�������G��d��U���u�u�u�%�g�<��������W9��h��U��%�e�4�%�6�<�(���B���F����ߊu�u�u�u�w�}�(߁�����R��[
�����2�i�u�
��1����	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��1����������^	�����0�&�u�x�w�}��������l��D�����2�
�'�6�m�-����
ۖ��l��_����4�%�4�%�2�q��������l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�g�<��������WO�C��U���u�u�u�u�w�-�G���	����]9��PN�U���
�9�=�n�w�}�W�������9F�N��U���u�
�
�9�?��������C9��V�����0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�H����l��A�����<�u�&�<�9�-����
���9F���*���
�%�#�1�>�����
����l��TN����0�&�%�d�:�%��������lW��V�����1�%�0�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����^��V�����u�=�;�_�w�}�W���Y�Ƽ�9��O1��*���
�;�&�2�k�}�(ށ�����l��d��U���u�0�&�u�w�}�W���Y����lW��V�����1�<�
�<�w�`��������C9��S1����u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�F�������@��V�����'�6�&�{�z�W�W���&¹��K9��h��*���<�;�%�:�w�}����
�μ�9��OB��*ۊ�4�
�'�2�w��(���&����_�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�4��-����PӒ��]FǻN��U���u�u�
�
�6��������C9��Z�����u�u�u�9�2�W�W���Y���F��1�����
�<�u�h�'�l����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�0�<�3�<�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�K����Z	��V�����;�&�2�4�$�:�(�������A	��D��*؊�0�<�1�4��1�[Ϯ�K����Z	��V�����'�2�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϮ�K����Z	��V�����u�=�;�_�w�}�W���Y�Ƽ�9��E��*���#�1�<�
�>�}�JϮ�K����Z	��V����u�u�u�u�2�.�W���Y���F���*���<�1�4�
�;��������C9��g�����%�#�1�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h>�����<�
�<�u�$�4�Ϯ�����F�=N��U���
�0�<�1�>�����
����l��TN����0�&�%�g��/���	�ԓ�V��S1�����%�g��'�8��������F��P��U���u�u�<�u��-��������Z��S��*؊�0�<�1�4��1�^������F�N��U���%�g��'�8��������C9��g����u�u�u�u�2�.�W���Y���F���*���<�1�<�
�>�}�JϮ�K����Z	��G��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠu�u�%�a��	����&����[��E��*ڊ�
�
� �d�f�<�(�������lǻN��Xʥ�a� ��8�9��(߁�	������^	�����0�&�u�x�w�}����,����Z��R1�����9�
�&�<�9�-����Y����V��V�����'�
�
�
�����H����W	��N��*���
�&�$���)�(���&��ƹF��R	�����u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�D������R��Y��]���6�;�!�9�0�>�G������lV��h\�� ��d�4�
�:�2�t�^Ϫ���ƹF�N��U���
�
�
�<�>�:��������WF������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�%�a��	����&����R��[
��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s�����h;�����2�0�d�i�w�/�(���&����U��_�����!�'�
�n�]�}�W��	�ғ�l2��^ �����4�
�9�u�$�4�Ϯ�����F�=N��U���
�
�<�<�0�8�F���&����R��P �����o�%�:�0�$�<�(���Y����U9��Q1�����f�
�%�1�9�q��������V��c1��F���8�g�_�u�w�8��ԜY���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��ي�&�
�|�4�3�3����	����@��X	��*���u�'�
�
���(���H�ד�C9��Y��\���=�;�_�u�w�}�W���Y����f9��Z��*���
�%�#�1�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����h;�����2�0�d�4��1�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(ځ�����C9��S1��*���u�&�<�;�'�2����Y��ƹF��h[�����4�
�9�
�9�.����
����C��T�����&�}�
�
�2�<��������lS��R�����9�
�'�2�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l��V1��*���|�u�=�;�]�}�W���Y���C9��U��*���#�1�<�
�>�}�JϮ�L����R9��h��N���u�u�u�0�$�}�W���Y���F��h[�����4�
�9�
�9�.���Y����Q��h�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W��	�ӓ�V��^ �����&�<�;�%�8�8����T�����h�����
�<�
�&�>�3����Y�Ƽ�\��DF��@���!�y�%�`�5�)�(����Ƽ�9��C�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`��������R��[
��U���;�_�u�u�w�}�W���&ƹ��G��Y1����u�
�
�0�6�W�W���Y�Ʃ�@�N��U���u�u�%�`�5�)�(���
���F��1�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�(ف�&����]��h^��Hʲ�%�3�e�3�e�;�(��&����V��Y1����u�x�u�
����������l��A�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��c�����
�
�%�#�3�<����&����\��E�����%�6�y�2�'�;�G���K����U��V�����u�%�&�2�4�8�(���
�Փ�@��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G�����:�}�4�
�8�.�(�������F��G1��E���g�3�
�f��-����P���G��d��U���u�u�u�%�a��#�������9��h��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}�(ف�&����]��h^�����1�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]ǑN�������8�;���W������lV��h\�� ��d�4�
�0�"�3�D�ԶY���F��1��!���;�
�
�
�'�+�Ͽ�
����C��R��U���u�u�%�c��	����&����R��[
�����;�%�:�u�w�/����Q����VJ��E��*ڊ�
�
� �d�f�<�(����ƭ�l��h�����
�!�
�&��t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�f�3�:�o�W���Y������T�����2�6�e�h�0�-�����ԓ�F9��1��*���0�|�|�!�2�}�W���Y���F��hX��*���<�2�0�d�6�����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�������8�;���(������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�}�WϮ�A����Z��P1��E��u�'�
�
���(���H�ד�C9��C��*��_�u�u�x�'�e� �������V9��V�����&�<�;�%�8�8����T�����h9�����2�0�e�4��1�(�������A	��N�����&�4�
�0�w�/�(���&����U��_�����;�y�4�
�>�����*���� 9��Z1����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GU��D��\ʴ�1�;�!�}�'�>��������lV�	��*���
�
�
� �f�l�������O��_�����u�u�u�u�w��(�������l��h�����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϮ�A����Z��P1��E���
�9�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���
�
�
�<�>�:���E�ƫ�C9��1��G���
�f�
�%�%�)����B���F���*���<�<�2�0�f�<�(���Y����T��E�����x�_�u�u���(�������lW��G1�����&�2�
�'�4�g��������C9��N�����e�3�g�3��n�(���������D�����
��&�f�1�0�E�ԜY�Ʈ�T��N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!��.�(�������\�V�����
�:�<�
�w�}����&ù��9��h_�*���1�;�|�|�w�5��ԜY���F�N��M���!�8�;�
���������R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�
�<�>�:��������WF������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����E]�