-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�_�&�w�8��������Z��X����_�0�!�!�w��5��=ǀ��l ��O��G���c�
�u�&�w�}�������9F�N��U���u�u�u�u�m�4�������W��N��U��������}�W�������	[�d��U���u�1�;�
��	�W�������AF��]����u�u�u�:�#�
�3���Cӏ��V��T��C�ߊu�u�n�u�w�-����s���F�S��U���;�u�!�
�8�4�(�������Z��`'��=��1�"�!�u�~�W�W���Y�ƨ�F���U���
�:�<�
�2�)�Ǻ�����w2��N�����u�|�u�u�~�W��������l��E����� �0�4�6�w�;����A�׈�U9��Q����;�
�a�d�>�W�W���T���K�C�X���x�x��8�8�8���T���K�C�X���x�_�u�u�8�-����Y����W����*���3�0�!�e�9�����Kӏ��F�N�����u�_�u�u�w�}�W���&����l��A�����u�u�u�;�w�)�(�����ƹF�N��U���
�-�&�4�#�<����Y�������*���<�
�0�!�%�n�W������]ǻN��U���u�u�
�-�$�/����&����Z���U���
�:�<�n�w�}�W���Y����l��D1�����
�1�!�u�m�2�ϭ�����Z��R����u�:�;�:�g�W�W���Y���9F���U���%�;�;�n�w�}�Z��T���K�C�X���u�:�4�u�>�3���T���K�C�X���u�u�&�2�6�}�(��������h����u�u�&�2�6�}�(��������h�����0�!�'�f�w�2����I��ƹF��^	��ʧ�!�4�<�u�w�)�(�����ƹF��^	��ʧ�!�4�4�u�w�)�(�������P��X����!�u�|�_�2�4�}���Y���K�C�X���x�x�x��$�<�������K�C�X���x�x�_�u�w��5��=ǀ��l��Q�����;�
�&�
�e�(�MϽ�����]��qV��Dۑ�3�e�4�
�'�%�(߁�����lU��N�����u�4�u�_�w�}�W���&����l��A�����u�u�k�4�#�<���Y���F��h�����!�4�4�u�w�}�J���&����RJǻN��U���
�-�&�'�$�1�(������F��C�����u�u�u�u�:�<��������l��C��H���
�1�!�_�w�}�L�ԜY���K�C�X���x�x�x�x��.�������K�C�X���x�x�x�_�w�}�(������F�UךU���
�1�!�u�k�}����&����{K��S�����u�k�r�r�w�5��������F�S��*����x�u�:�9�2�G��YԾ�F��EN����h�}�1�;���#��Y����G	�S�R��|�u�9�0�3�3�L���Yӂ��GF�N�U���1�!�n�_�9�}��������A��