-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�m�m�d�a���(���
����GF�N�����9�u�u����;���:���F��h��U���������}���Y����G��T��;ʆ�����]�}�W�������	F��cN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�%�<���6����g"��x)��N���u�<�
�9�?��W���7ӵ��l*��~-��0����}�d�1� �)�W���s���Z��V��U���������!���6���F��@ ��U���_�u�u�;�5�)�(���Y����g"��x)��*�����}�d�3�*����P���F��h�� ���e�o�����;���:����g)��]����!�u�|�_�w�}��������F��x;��&���������W��Y����G	�UךU���%�'�!�'��}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y����C9��C��*���u� �u����>���<����N��S�����|�_�u�u�'�>�W���7ӵ��l*��~-��N��1�_�_�'�?�)����ӄ��R��QN��M��d�a�
�
��}��ԜY�Ư�]��Y�����;�!�9�2�4�l�Mύ�=����z%�
N��R�ߊu�u�:�&�6�)��������_	��T1�Oʆ�����m�}�G��Y����\��V ������&�d�3�:�m�Mύ�=����z%��r-��'���e�1�"�!�w�t�M���I����V��^�E��e�e�w�_�w�}��������C9��h��*���
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��_�N���u�6�;�!�9�}����&����U��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��H���9F������!�4�
��$�i����J����g"��x)��*�����}�e�3�*����P���V��^�E��e�e�e�d�g��}���Y����G����&���!�
�&�
�w�}�#���6����e#��x<��G���:�;�:�e�w�`�U��I����V��^�D��e�n�u�u�4�3����Y����g9��1�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��UךU���:�&�4�!�6��#���N����lP�=��*����
����u�GϺ�����O�
N��E��e�e�e�e�g�m�G��[���F��Y�����%��
�!��.�(���Y����)��t1��6���u�g�u�:�9�2�G���D����V��^�E��e�e�e�e�l�}�WϽ�����GF��h=�����3�8�m�o���;���:����g)��\����!�u�|�o�w�m�G��I����W��^�E���_�u�u�:�$�<�Ͽ�&����GW��Q��L��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��	���&����V�=��*����
����u�GϺ�����O�
N��E��e�e�e�e�g�m�G��[���F��Y�����%��
�!�e�;���Y�Ɵ�w9��p'��#����u�g�u�8�3���Y���V��^�E��e�e�e�e�g�f�W�������R��V��!���d�
�&�
�e�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����W��^�E��e�w�_�u�w�2����Ӈ��`2��C_�����d�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�N���u�6�;�!�9�}����&����l ��h_�Oʆ�������8���K�ƨ�D��^��O���e�e�e�d�g�m�G��I����]ǻN�����4�!�4�
��.�Fف�
����\��c*��:���
�����m��������\�^�E��e�e�e�e�g�m�G���s���P	��C��U����
�!�b�1�0�F���Y����)��t1��6���u�g�u�:�9�2�G���D����V��^�E��e�e�e�e�l�}�WϽ�����GF��h=����
�&�
�b�m��3���>����v%��eN��Eʱ�"�!�u�|�m�}�G��I����V��^�E��w�_�u�u�8�.��������l��1����u�u��
���(���-���V��X����u�h�w�e�g�m�G��I����V��L�U���6�;�!�;�w�-�$����֓�@��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I���9F������!�4�
��$�o�(���&���5��h"��<������}�g�9� ���Y���F�^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���P	��C��U���6�;�!�9�f�l�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��H����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����W��d��Uʶ�;�!�;�u�'�>��������T�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����W��^�����u�:�&�4�#�<�(���
���� T��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��h\��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�D���_�u�u�:�$�<�Ͽ�&����G9��\��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[�*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��F؊�f�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��d�e�d�n�w�}��������R��X ��*���g�f�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�d�l�}�WϽ�����GF��h�����#�g�l�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�f�f�W�������R��V�����
�#�g��m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�f�l�L���YӅ��@��CN��*���&�
�#�g�f�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���P	��C��U���6�;�!�9�d��1���<���5��h"��<������}�f�9� ���Y���F�_�D��e�d�e�d�f�m�F��I����V�=N��U���&�4�!�4��2�����ԓ�u^��^�Oʆ�������8���J�ƨ�D��^��O���e�d�d�d�f�m�G��I����V��^�E��n�u�u�6�9�)����	����@��A]��D���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��F؊�b�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��d�d�d�n�w�}��������R��X ��*���g�d�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�d�d�u�W�W�������]��G1�����9�m��u�w�	�(���0����p2��F����!�u�|�o�w�l�F��H����F�T�����u�%�6�;�#�1�E܁�Y�Ɵ�w9��p'��#����u�g�u�8�3���Y���V��^�E��e�e�e�e�g�m�L���YӅ��@��CN��*���&�
�#�g�o�m�G��Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)����I����g"��x)��*�����}�u�8�3���Y���V�=N��U���&�4�!�4��2��������	F��s1��2������u�e�9� ���Y���F�_�����u�:�&�4�#�<�(���
���� 9��N��1��������}�EϺ�����O�
N��D���_�u�u�:�$�<�Ͽ�&����G9��1�Oʆ�������8���Kӂ��]��G��H���d�w�_�u�w�2����Ӈ��P	��C1��F��o������!���6�����Y��E���h�w�e�w�]�}�W���
������T�����f�f�o����0���/����aF�
�����e�u�h�w�f��}���Y����G�������!�9�f�g�m��3���>����v%��eN��U���;�:�e�u�j��F���s���P	��C��U���6�;�!�9�d�i�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���I����F�T�����u�%�6�;�#�1�O��Cӵ��l*��~-��0����}�u�:�9�2�G���D����V��^�����u�:�&�4�#�<�(���
����S��^�Oʆ�������8���H�ƨ�D��^��O���d�e�e�e�g�m�G��B�����D��ʴ�
�:�&�
�!�h�C��Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�n�u�w�>�����ƭ�l��D�����`�e�o����0���/����aF�N�����u�|�o�u�g�m�F��I����V�=N��U���&�4�!�4��2�����ӓ�V�=��*����
����u�CϺ�����O�
N��E��e�e�e�e�g��}���Y����G�������!�9�d�
�g�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��u�u�6�;�#�3�W�������l
��1�Oʆ�������8���K�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-��������9��q(��3���o������!���6��� F��@ ��U���o�u�d�d�f�l�F��H����W��_�D��d�d�d�n�w�}��������R��X ��*���a��u�u���8���&����|4�]�����:�e�u�h�u�m�G��I����V��^�E��e�d�d�d�f��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�m�G���s���P	��C��U���6�;�!�9�d��1��I���5��h"��<������}�f�9� ���Y���F�_�D��d�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��2��������	F��s1��2������u�f�9� ���Y���F�L�U���6�;�!�;�w�-��������9��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}��������ES��T��!�����
����_�������V�S��E��e�n�u�u�4�3����Y����\��h��*���u��
����2���+����W	��C��\��u�e�e�d�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�g�l�G��Y����\��V �����:�&�
�#��}�W���&����p9��t:��U��1�"�!�u�~�g�W��B���F��P ��U����
�&�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��n�u�u�4�#�4��������]��^ ��Oʦ�'�;�n�u�w�<��������@��Y�����:�u�%���.�W��������� ����u�u�&�2�6�}��������B9��h��*���
�u�u����>��Y����Z��[N��*���
�1�
�l�m��8���7���F��P ��U���
� �l�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h_�U����
�����#���Q����\��XN�N���u�&�2�4�w�-��������`2��CX�����u�u��
���L���Yӕ��]��V�����1�
�d�o���2���s���@��V�����2�6�0�
��.�Fف�
����\��c*��:���n�u�u�&�0�<�W���
����W��N�7�����_�u�w�4��������S�=��*����
����u�FϺ�����O��N�����4�u�%�&�0�>����-����l ��hV��U���
���n�w�}�����ƭ�l��h��*��o�����W�W���������D�����
��&�d��.�(��Cӵ��l*��~-�U���&�2�4�u�'�.��������	F��x"��;�ߊu�u�<�;�;�<�(���&����l5��D�*���
�m�o����0���s���@��V�����2�7�1�l�w�}�8���8��ƹF��^	��ʳ�
��-� ��k�(���H�ޓ�F��d:��9�������w�n�W������]ǻN�����9�3�
��/�(�(��&����U��T��!�����
����_������\F��d��Uʦ�2�4�u�%�$�:����&����GT��D��U����
���l�}�Wϭ�����R��^	�����d�u�u����L���Yӕ��]��C��G���
�e�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��E��D��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����;����G9�� 1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������`��C1�B���2�d�f�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��G���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����A��]�U����
�����#���Q�ƨ�D��^����u�<�;�9�1��5�������
9��Q��CҊ�d�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�&����|��X��G���2�d�`�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ʈ�\
��p+�� ���c�
� �f�o�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��X������!�d�a�%�:�F��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����
� �a�f�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h�����f�f�o����0���/����aF�
�����e�n�u�u�$�:����	����l��F1��*���
�&�
�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�1��n�W���6����}]ǻN�����9�3�
�!�n��(���L�ѓ� F��d:��9�������w�n�W������]ǻN�����9�3�
�!�n��(���&����\��c*��:���
�����l��������l�N�����u��6�
�e��(���L�ғ� F��d:��9�������w�n�W������]ǻN�����9�3�
�!�f�m�B�������F��d:��9�������w�n�W������]ǻN�����9�3�
�!�f�n�C���&����CU�=��*����
����u�FϺ�����O��N�����4�u��6��l�(ہ�����
V�=��*����
����u�FϺ�����O��N�����4�u��6��o�(ہ�����l��N��1��������}�D�������V�=N��U���;�9�3�
�#�l�G������� _��N��1��������}�D�������V�=N��U���;�9�:�!��>����J����G��D�����
�`�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƣ�G9��T��*���"�<�0�4�$�:�(���&����\��c*��:���
�����}�������9F������:�
�:�1��i����Aù��\��c*��:���
�����}�������9F������:�
�:�1��i����H����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�d��(�@���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�d�
�2��C��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�b�3�
�e��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����b�'�2�d�f�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��Dӊ� �b�l�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���
�a�c�o���;���:����g)��^�����:�e�n�u�w�.����Y����U��]��G��������4���Y����W	��C��\�ߊu�u�<�;�;�;�(���=����lW��h��*��f�o�����4���:����U��S�����|�_�u�u�>�3�Ͽ�&����P��h=�����3�8�c�o���;���:���F��P ��U���&�2�7�1�f�i�MϜ�6����l�N�����u��-� ��3����Nƹ��U��Y��F��������4���Y����W	��C��\�ߊu�u�<�;�;�;�(���5�Ԣ�F�� [��*���
�a�f�o���;���:����g)��]����!�u�|�_�w�}����Ӈ��@��T��*���&�d�
�&��o�Mύ�=����z%��N�����4�u�%�&�0�?���M����|)��v �U���&�2�4�u��>�(�������F��E��G���3�
�b�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W������� ��T������'�6� �2�i�(ց�����R�=��*����
����u�FϺ�����O��N�����4�u�%�&�0�>����-����9��Z1�U����
���l�}�Wϭ�����R��^	�����m�u�u����L���Yӕ��]��Q=�����&�
�!� �#�/�(���@����V��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�1�����
����A��B��Aӊ�
�0�
�a�g�g�$���5����l0��c!��]��1�"�!�u�~�W�W������� ��T������'�6� �2�h�(ׁ�����
9��T��!�����
����_������\F��d��Uʦ�2�4�u��4�����*����G��h[��M���2�d�c�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h
�����;�3�
�e�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��B���8�'�4�
�2��C��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
� �d�m��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���
�a�b�o���;���:����g)��^�����:�e�n�u�w�.����Y����G��_�����2�;�3�
�g�o����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���d�d�1�8�%�<�(���&����\��c*��:���
�����}�������9F������!�%�g�
�2�2��������^��N�&���������W������\F��d��Uʦ�2�4�u�8��h��������A��Z�U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Dׁ�����9��T��!�����
����_�������V�=N��U���;�9�!�%�d�����M���5��h"��<������}�w�2����I��ƹF��^	��ʦ�9�!�%�e��8��������W��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����H����\��Y1����l�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����W��E	��*���d�m�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��h
�����;�'�2�d�g�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������hZ�����g�b�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lR��E��D��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������9��Z����� �d�d�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��Dۊ�0�:�2�;�%�:�F��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V����� �l�
�e�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��B1�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������V��c1��A���8�f�o����0���s���@��V�����2�7�1�g�`�g�5���<����F�D�����%�&�2�6�2��#���Hù��^9��N��1�����_�u�w�4��������T9��S1�A������]�}�W�������C9��P1������&�d�
�$��D��*����|!��d��Uʦ�2�4�u�%�$�:����K���$��{+��N���u�&�2�4�w�-��������`2��C_�����d�u�u����>��Y����Z��[N��*���
�1�
�f�w�}�8���8��ƹF��^	��ʲ�%�3�
�e��m�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�� ��f�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����q5��B��Cӊ� �d�m�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����U5��u=�� ���c�
� �d�o�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����d�
�e�o���;���:����g)��]����!�u�|�_�w�}����Ӂ��l ��_�����u��
����2���+������Y��E��u�u�&�2�6�}��������B9��h��D���8�g�u�u���8���B�����Y�����<�
�1�
�b�}�W���5����9F������2�%�3�
�e��G��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��	��*���d�e�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��h_�*��o������!���6���F��@ ��U���_�u�u�<�9�1����;����G9��Q��D݊�f�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����T��G_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u���$�������lW��B1�G���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&���� R��N�&���������W������\F��d��Uʦ�2�4�u�'��(�F���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
� �d�l�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��D���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϲ�	����R��G^��U���
���
��	�%���Y����G	�UךU���<�;�9�2�'�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʲ�%�3�
�`��m�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������[��h�����3�
�b�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��D���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	�ד�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�2��������9��T��!�����
����_�������V�=N��U���;�9�;�!�?����A����	F��s1��2������u�g�9� ���Y����F�D���������#�l�@�������V��G\��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%����M����	F��s1��2������u�g�9� ���Y����F�D���������#�l�N�������G9��h\�*��o������!���6���F��@ ��U���_�u�u�<�9�1����Hù��lT��h�Oʆ�������8���Nӂ��]��G�U���&�2�4�u�:��D���&����CW�=��*����
����u�EϺ�����O��N�����4�u�:�'�$����@����	F��s1��2������u�g�9� ���Y����F�D�����:�9�&�
�"�o�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V��&�����!�d�n�3����&����CT�=��*����
����u�FϺ�����O��N�����4�u�'�
�"�l�N���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V��&�����!�!��3�(���K�֓�F��d:��9�������w�n�W������]ǻN�����9�3�
��/�(�(݁�����l ��W�����u��
����2���+������Y��E��u�u�&�2�6�}����@����^��GZ��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�o�(���K�ғ�F��d:��9�������w�o�W������]ǻN�����9�;�!�=�c�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʻ�!�=�a�3��l�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
� �f�g�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h\�����d�
�d�o���;���:����g)��\����!�u�|�_�w�}����ӈ��A��h��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϰ�����l ��]�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����^��N�&���������W������\F��d��Uʦ�2�4�u�8��i����MŹ��\��c*��:���
�����}�������9F������!�%�g�
�"�n�E���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����b�3�
�b��n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���f�a�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӏ��C9��h]�*��o������!���6�����Y��E��u�u�&�2�6�}��������l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�l����Hƹ��\��c*��:���
�����}�������9F������&�9�!�%��(�C���	����`2��{!��6�����u�e�3�*����P���F��P ��U���6�
�l�d�1��Gց�J����g"��x)��*�����}�d�3�*����P���F��P ��U���%�;�!�3��i�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����3�
�l�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��*���a�c�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l�� 1��*���
�g�o����0���/����aF�
�����e�n�u�u�$�:����*����
_��h��A���%�u�u����>���<����N��
�����e�n�u�u�$�:��������CP��R�����3�
�f�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��F���8�'�4�
�"�i�C���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����
� �f�b�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��*���a�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:����*����
_��h��A���%�u�u����>���<����N��
�����e�n�u�u�$�:��������CT��S�����
� �a�l�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��@���
�l�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��GV�� ���d�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������l_��1��*��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������lW��h��@���%�u�u����>���<����N��
�����e�n�u�u�$�:����*����T��1��*��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������lW��h]�� ���b�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G9��1��*��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������lW��h\�� ���b�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G9��1�����`�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӏ��P��]��*���`�d�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�l��\��C���
�b�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������`9��h_�*݊� �`�d�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����U5��C1�E���3�
�m�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W������� ��T��Gڊ�
� �`�`�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h�����
�d�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƣ�D5��h�����&�
� �c�n�-�W���-����t/��a+��:���g�1�"�!�w�t�}���Y����R
��R�����
�g�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƣ�l��S_�� ��d�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������]��Q��@ي�g�o�����4���:����V��X����n�u�u�&�0�<�W���*����U��[��F��������4���Y����\��XN�N���u�&�2�4�w�8�$���&���� Q��N�&���������W������\F��d��Uʦ�2�4�u�8��o����OĹ��\��c*��:���
�����}�������9F������<�8�b�3��j�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����;�!�3�
�n��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��D؊� �c�c�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���c�m�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��Z�����'�4�
� �`�d����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���d�
� �b�b�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����m�1�8�'�6����N����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�d��(�@���	����`2��{!��6�����u�e�3�*����P���F��P ��U���-��,� ��9�(��&����S��N�&���������W��Y����G	�UךU���<�;�9�9�4�����Mʹ��\��c*��:���
�����}�������9F������9�6��d�1��Bց�H����g"��x)��*�����}�g�3�*����P���F��P ��U���
�
�
�f�1��Aց�K����g"��x)��*�����}�u�8�3���B�����Y�����<�<�3�
�a��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��E�����3�
�b�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������hY�����3�
�m�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��*���m�`�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��^�� ��d�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������l��h�����&�
� �b�n�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��D�����
� �b�b�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��e�����
� �m�`�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��9����!�d�`�>�����&¹��l^��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�#�-�D���&����CT�=��*����
����u�W������]ǻN�����9�!�%�`�1��Cځ�K����g"��x)��*�����}�u�8�3���B�����Y�����g�
� �m�f�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��L���
�c�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��h��M���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����U�� Y��F��������4���Y����\��XN�N���u�&�2�4�w��F���H����S��G]��U���
���
��	�%���Kӂ��]��G�U���&�2�4�u�:��@���&����CU�=��*����
����u�GϺ�����O��N�����4�u�
�0�"�)�Fށ�����l��N��1��������}�D�������V�=N��U���;�9�3�
���E�������l��Q����� �m�b�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����@��C��D���
�e�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G_�����d�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����G��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:����*����2��x��D���3�
�e�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W������� ��T������'�6� �2�i�(݁�����l��N��1��������}�D�������V�=N��U���;�9�3�
�#���������F��\�� ��a�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G9��D�����!�'�
�g�c�;�(��&���5��h"��<������}�f�9� ���Y����F�D������6�
�4�2���������9��Q��C݊�f�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�&����R��d�����0�a�
� �n�l����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*����&�
�!�"�)����@�ד�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w���������G��C��*���g�3�
�m��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��d1��*���0��'�6�"�8�Cց�&����
S��N�&���������W��Y����G	�UךU���<�;�9�3��)�4���&����P��R1�*���l�m�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�l��t��*��� �!�'�
�a�l����I�ߓ� F��d:��9�������w�n�W������]ǻN�����9�3�
�!��.�(�������V9��h\�� ��d�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӏ��P��V��&���6� �0�`�����K����\��c*��:���
�����l��������l�N�����u�
�4�g�f�;�(��N����	F��s1��2������u�d�}�������9F������9�6��g�1��G���	����`2��{!��6�����u�b�3�*����P���F��P ��U���
�
�
� �f�h�(��Cӵ��l*��~-��0����}�g�1� �)�W���s���@��V�����
�d�3�
�g�h����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���d�d�
� �f�k�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����c�3�
�e�n�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��X��܊� �d�b�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����T��Q��Aފ�g�o�����4���:����V��X����n�u�u�&�0�<�W����ԓ�l ��^�*��o������!���6���F��@ ��U���_�u�u�<�9�1����/�ғ�F9��\��A��������4���Y����\��XN�N���u�&�2�4�w�2�(���&����W��G_��U���
���
��	�%���Kӂ��]��G�U���&�2�4�u�:��(�������P��N�&���������W������\F��d��Uʦ�2�4�u�8���C��&����T��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�;�#�5�O���&����l��N��1��������}�GϺ�����O��N�����4�u�:�9�$����Jǹ��\��c*��:���
�����}�������9F������2�%�3�
�c��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��G1��؊�
� �d�`��l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��X��*܊� �d�c�
�c�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����_	��a1�����d�f�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��^Y�� ��b�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����Z9��h_�����d�f�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӈ��A��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������9��h_�@���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�G���&����l��N��1��������}�D�������V�=N��U���;�9�3�
�2�0�(���+����l��h-�����b�3�
�g�d�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��D�����d�3�
�g�f�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��Q=�����
�;��;�2�<��������9��h_�A���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����9��h_�G���u�u��
���(���-��� W��X����n�u�u�&�0�<�W�������l/��e�����1��0�6���(���H����CU�=��*����
����u�FϺ�����O��N�����4�u� �
�'�/����J����G��D�����
�g�l�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����\��a�����
�
�'�!��.��������^��N�&���������W��Y����G	�UךU���<�;�9�:�#�
��������D��R1�����
� �d�f��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��R����
�4�!�3��o�G���Y�Ɵ�w9��p'��#����u�b�1� �)�W���s���@��V����� �l�
�%�8�8�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1��*���6�u�u����>��Y����Z��[N��*���
�&�$���)�(���&����`2��{!��6�ߊu�u�<�;�;�<�(���&����
V��N��:����_�u�u�>�3�Ϲ�	����V��T��U���
���n�w�}�����ƫ�C9��h_�*���:�0�o����0���/����aF�
�����e�n�u�u�$�:��������lW��h�����o������!���6�����Y��E��u�u�&�2�6�}��������l	��X
��Oʆ�������8���Mӂ��]��G�U���&�2�4�u�'��(���Y�Ɵ�w9��p'��#����u�g�u�8�3���B���F��Z�����8�m�m�d�c��(�������lU��D1����g�f�3�9��.�W���Y����V��^�����u�u�u��m��#���+���F�N��8�����o����%�ԜY���F��Y^��<���u�u����f�W���Y����Z��`'��=������]�}�W���Y����l1��c&��U�����u�n�w�}����Y���F�N�����u��
���L���Y�����R��U��������W�W���Y�ƨ�]V�'��&���������W��Y����G	�UךU���u�u�<�d�m��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����C��RN�<����
�����#���Q�ƨ�D��^����u�u�u�0�m��W���&����p]ǻN��U���:�!�o����3���>����v%��eN��Dʱ�"�!�u�|�~�W�W����Ư�^��R ���ߊu�u�:�%�9�3�W���;���� ��h����;�
�g�&�d��(�������/��N�����'�6�}�u�w�}�Wϗ�Y�ƅ�g#��eUךU���u�u� �
���W���7����a]ǻN��U���<�e����g�>���>����F�N�����
���u�w��2���B���F�
�������o����%���s���C	��FךU���u�u�9�u�w��$���5����l�N��Uʧ�&�!�o��w�	�(���0��ƹF�N����o��u����>���<����N��
�����e�n�u�u�w�}����Y�ƅ�5��h"��<������}�f�9� ���Y����F�N�����u������4�ԜY���F��B��U���u��
����2���+������Y��E���n�u�u�0�3�>��������9l�N�����0�!�8�m�o�l�C���&����lU��D1����g�d�8�-�3�-�>�ԜY�ƫ�]��TN��U���u�u��u�w��2���B���F� ��*����u�u����L���Y�����1��1���o�����W�W���Y�ƨ�]W��~*��U������n�w�}�W�������d/��N�<�����|�_�w�}����Q���F�
��E���u��
���(���-��� W��X����n�u�u�u�w�9����Y����g"��x)��*�����}�d�3�*����P���F�N�� ���u� �u����>���<����N��
�����e�u�n�u�w�8�Ͻ�����]��=d��Uʶ�8�:�0�!�:�e�O���M����U��h]����;�
�
�u��}�WϹ�����NǻN��U����o�����}���Y���}3��d:��0������]�}�W���Y����l1��c&��U�����n�u�w�}�WϺ�¹��w2��N��!����_�u�u�w�}����.����\��y:��0���n�u�u�%�%�}�}���Y���W��T��;ʆ�������8���J�ƨ�D��^����u�u�u�<�f�g�>���-����t/��a+��:���f�u�:�;�8�m�L���Y���	��X
��Oʜ�u��
����2���+����W	��C��\�ߊu�u�u�u�8�)�Mϑ�-ӵ��l*��~-��0����}�u�:�9�2�G���B����������;�n�_�_�2�4�}���Y����U��Q��*���&�f�;�
�e�n����&����fV������;�u���f���������@��\��*���&�f�
�
�"�1����Y����V��^�����_�u�u�u�w��J���U���F� ��*����u�k�f�]�}�W���Y����l1��c&��K��y�u�u�u�w�9�ށ�0����X�BךU���u�u�:�!� ��?��Y���F�G��U���u�_�u�u�w�}����GӇ��P
��=N��U���u�0�0�u�i�<�(���U���F�
��E��u�'�
� �n��G�ԜY���F��Y_��Kʲ�%�3�
�l�'�q�W���Y����C��RN��U���
� �l�
�'�2��ԜY���F��S����3�
�l�6�{�}�W���Yӂ��GF�	��*���l�
�g�n�]�}�W���&����lU��D1����g�f�3�9��.�(��CӅ��C	��Y��3җ�d��3�e�1�9�(���
����@9��h]�� ���1�%�u�u�0�3�������9F�N��U���h�u�y�u�w�}�Wϐ�4����t#�	N����u�u�u�<�g�
�3���D����l�N��Uʱ�;�
���w�c�D��Y���F��X��"����h�u�g�]�}�W���Ӌ��NǻN��U���9�u�k�4��1�[���Y�����R��Kʴ�
�&�y�u�w�}�WϺ������h��D���%�y�u�u�w�}����Y����A��B1�F���y�u�u�u�w�>�W�������F9��1��Y���u�u�u�1�"�}�IϹ�	����V��G\����u�3�e�3�"��E���J���� T��h��*���
�g�o�6�:�2�����ގ�W��Q1�����
�g�&�f�9��E�������@ǻN�����<�u�4�u�]�}�W���Y���F��=N��U���u� �
���}�I��s���F�S��*����u�k�f�{�}�W���Yӂ��9��s:��H���g�_�u�u�w�}����.����[�\��U���%�'�u�4�w�W�W���Y�ƨ�]V�	N��*���-� �
�c��(�F���	��ƹF�N����h�u�������@����V��G_�U���u�u�1� �w�c����;����G9��1��*��
�g�n�_�w�}�(߁�������\��*ۊ�
�f�o�6�:�2�����ގ�W��Q1�����
�g�&�f�9��(�ԜY�ƫ�]��TN�����u�u�u�u��}�I��s���F�y;��&����h�u�y�w�}�W�������d/��N��U��_�u�u�u�w�4�F���=���F��d��U���u�1� �
��	�W���H���F��E�����_�u�u�u�w�4�G��Y����U��Z��E�ߊu�u�u�u�>�l�J�������lW��h����u�u�u�%�8�8�J�������lW��h�����_�u�u�u�w�2���Y����U��Z��G��_�u�u�
��>�������]��h_��A��6�8�:�0�#�0�O��H�Ҫ�9��Z��G���f�;�
�
�]�}�W�������^��d��U���u��u�k�f�W�W���Y�Ƃ�~9��v)��H���y�u�u�u�w�9�߁�0����X�BךU���u�u�<�d� ��?��Y����F�N�����
���u�i�l�}���Y������FךU���u�u�<�e�j�}��������l��=N��U���u�<�d�h�w�/�(���H�֓�JǻN��U���%�:�0�h�w�/�(���H�֓�C��RBךU���u�u�:�!�j�}��������l��dךU���
�
�6�%�d�3�(���
�ד�l3��N�����0�!�8�m�o�l�C���&����lU��D1����
�_�u�u�2�8�������F�N��<���k�d�_�u�w�}�W���&����vF�_�U���u�u�1�;���#���G����9F�N��U���d����j�}�E�ԜY���F��B��<���u�k�d�_�w�}�������9F�N��U���e�h�u�'��(�F���	��ƹF�N����h�u�'�
�"�l�B���U���F������h�u�'�
�"�l�B�������9F�N��U���!�h�u�'��(�F���	����9lǑ=N��U���!�0�6�'�2�)�����έ�l%��Q��U���!�0�&�4�2�0�������9F���6���&�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�}���Y���F�N��U���4�
��3�:�a�W���7����^]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p�����Ƽ�\��D@��X���u�%�:�0�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�d�|�!�2�W�W���Y���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��؊�&�
�|�|�#�8�}���Y���F�N�����
��,� ��k�(���&����Z�U��*���,� �
�c��(�D���	��ƹF�N��U���u�u�������N����lW��N�U������!�f�j����H����l�N��U���u�u�u�3������&����9��P1�@���h�3�
��/�(�(��&����lT��h����u�u�u�u�w�}�W���&�ғ�V��Z�I���8�
�a�3��h�(��s���F�N��U���!�%�g�'�0�l�D���DӒ��lT��B1�E���n�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9l�N�U���<�;�%�:�2�.�W��Y����A	��D�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���O��_��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����VO��Y
�����4�
�!�'�w�}��������\��h^��\���=�;�u�u�w�}�W���Y����`9��d����l�'�2�d�f�}�Jϸ�&����|��X�����e�
�g�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dךU���x�4�&�2�w�/����W���F�G�����}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�I�����_�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��h\��\ʡ�0�_�u�u�w�}�W���Y�ƪ�l��_��A���2�d�l�u�j�;�(���H�Փ�l ��X����u�u�u�u�w�}�W�������lW��hZ�����f�`�i�u��>�(��&ǹ��lP��h����u�u�u�u�w�}�W�������9��E��D��u�h�3�
�#�l�G�������9��d��U���u�u�u�u�w�;�(���@ʹ��A��]�U��3�
�!�l�����N����9F�N��U���u�u�u�'�4�3�F��&����R��R�����:�1�
�a�1��O߁�K���F�N��U���u�:�!��4�2�(�������l��^	�����d�e�u�h�8�)�$�������l��C�����;�3�
�`��n�}���Y���F�N�����!�%�`�'�0�l�F���Dӕ��l��[�� ��f�%�n�u�w�}�W���Y�����h��D݊�0�
�a�l�k�}��������U��_��G�ߊu�u�u�u�w�}�W�������CW��E��D��u�h�&�9�#�-�N���&����CT��N��U���u�u�u�u�#�-�������� F���*��� �a�f�%�l�}�W���Y����������u�u�u�;�w�;�}���Y����C��R�����u�x�u�&�>�3�������KǻN�����&�u�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��R���=�;�u�u�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��|�u�=�;�w�}�W���Y���F��d1��*���0��'�6�"�8�C݁�&����R��R�����!��&�
�#�(����&�ԓ�l ��Y����u�u�u�u�w�}�W�������l%��R1����� �0�a�
��8�(��I���U5��C1�����!� �!�'��d�N���&����l��=N��U���u�u�u�u�w���������G��C��*���m�'�2�d�a�}�Jϸ�&����R��d�����0�`�
�
�"�l�Eց�J���F�N��U���u�&�9�!�'�d�(�������l��h_�G��u�0�
�8�f�l��������U��W����u�u�u�u�w�}�W���
����^��1�����4�
�0�
�c�j�K�������CT��h
�����;�3�
�d�d�-�L���Y���F�N��U���
�8�g�d�3�0����&����S��R�����!�%�d�
�2�2��������R��UךU���u�u�u�u�w�}����N����\��Y1����b�u�h�!�'�l�(�������l ��^�*��_�u�u�u�w�}�W���Y����S��R�����'�2�d�m�w�`����Kƹ��^	��V �� ��g�
�g�_�w�}�W���Y���F��G1�*���:�2�;�'�0�l�G���DӒ��lU��S�����
� �d�m��o�}���Y���F�N�����f�
�0�
�c�j�K�������l ��^�*��_�u�u�u�w�}�W���Y���� ^��R	��A��i�u�8�
�o�;�(��O����9F�N��U���u�u�u�8��n����H����[��Z��F���
�g�b�%�l�}�W���Y����������u�u�u�;�w�;�}���Y����C��R�����u�x�u�&�>�3�������KǻN�����&�u�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��R���=�;�u�u�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��Q��@���u�=�;�u�w�}�W���Y��� ��O/�����
�m�
�0��i�D��Y����U��]��G�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�F܁�
����O�C�����u�u�u�u�w�}�W���������C1�@���'�2�d�a�w�`����4����])��h_�*ي� �l�b�%�l�}�W���Y����������u�u�u�;�w�;�}���Y����C��R�����u�x�u�&�>�3�������KǻN�����&�u�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��R���=�;�u�u�w�}�W������N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��h��*���u�'�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�a�;���P���G��=N��U���u�u�u�u�w�8�(��Y����A��B1�*��_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9F�C����2�u�'�6�$�s�Z�ԜY�Ƽ�\��DN�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D����F��R ךU���u�u�u�u�1�u�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O�X��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�d�~�2�W���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���Hʹ��^9��G��U���;�u�u�u�w�}�W���YӔ��lW��R�����3�
�l�%�l�}�W���Y����������u�u�u�;�w�;�}���Y����C��R�����u�x�u�=�w�8�ϭ����R��d1�����3�!�0�&�6�8�������KǻN�����
�&�
�&�>�3����Y�Ƽ�\��DN�����4�!�u�%���������l�N�����u�u�u�u�4�.�W���:����^F��=N��U���u�u�u�=�9�<�(���
�ד�@��S����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t�������R��C��U���%�6�;�!�;�:���P����[��N��U���u�u�u�u�w�}����*����Z�V��!���g�3�8�d�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:��؊�&�
�u�k�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W�������l ��R������&�f�3�:�o�}���Y���F�N�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�����B���F�N��U���u�;�u�3�]�}�W���Y���D����&���!�
�&�
�w�c�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�c�;���s���F�N��U���0�&�_�u�w�}�W���Y���F�V��&���8�i�u�%���܁�
����9F�N��U���u�u�u�;�w�;�}���Y���F�@��U����
�!�
�$��W���s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�B�������F�N��U���u�u�0�&�]�}�W���Y���F�N������3�8�i�w�-�$���ǹ��^9��=N��U���u�u�u�u�w�3�W���s���F�N�����u�%��
�#�����Y���F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����
�&�u�h�6��#���O����lS��N��U���u�u�u�u�2�.�}���Y���F�N��U���4�
��3�:�a�W���*����9��Z1����u�u�u�u�w�}�W���Y����F�N��U���"�0�u�%���ف�
����X�N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���%��
�&�w�`����-����l ��hX�U���u�u�u�u�w�}����s���F�N��U���u�u�4�
��;���Y����g9��1�����_�u�u�u�w�}�W���Y����Z ��N��U���u�u�"�0�w�-�$���Ĺ��^9��
P��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}�W�������F�N��U���u�u�u�u�6��$������R��c1��B���8�c�_�u�w�}�W���Y���V��^�U���u�u�u�u� �8�W���*����9��Z1�H���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W���Y����_��N��U���u�u�u�u�w�}����*����Z�V��!���m�3�8�b�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����g9��1����h�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���e�3�8�l�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:�����3�8�l�h�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�d�1�0�F��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�F߁�
����9F�N��U���u�u�u�;�w�;�}���Y���F�@��U����
�!�d�1�0�F���G���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���;���&�u�h�4��	���&����W��N��U���u�u�u�u�2�.�}���Y���F�N��U���4�
��3�:�a�W���*����W��D��E�ߊu�u�u�u�w�}�W����ƥ�l�N��U���u�"�0�u�'��(���K����lW��
P��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�%���.�W������l��1����n�u�u�u�w�}�W���YӃ��Vl�N��U���u�u�u�u�w�<�(������F��h=����
�&�
�d�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����g9��]�����g�h�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���7����^F���&���!�a�3�8�f�f�W���Y���F�N�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�f�����K���F�N��U���u�0�1�<�l�}�W���Y�����YN��*���&�d�
�&��n�J���Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��h �����i�u�%���)�B�������9F�N��U���u�u�u�9�2�}�W���Y���F�N��U����
�&�u�j�<�(���
����U��]�U���u�u�u�u�w�}������ƹF�N��U���=�;�4�
��.�Fځ�
����[�=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���4�
��3�:�a�W���*����P��D��@�ߊu�u�u�u�w�}�W�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��@���8�d�n�u�w�}�W���Y����������u�u�u�u�w�5�Ͽ�&����GW��Q��D���k�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�<�(������F��h=����
�&�
�c�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�c�1�0�F��Y���F�N��U���;�u�3�_�w�}�W���Y�ƻ�V��G1��*���b�3�8�d�w�c�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�f�����N���F�N��U���u�0�&�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���N����lW��=N��U���u�u�u�u�w�3�W���s���F�N�����u�%��
�#�e����H���l�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U����
�&�u�j�<�(���
����U��V�U���u�u�u�u�w�}����s���F�N��U���u�u�4�
��;���Y����g9��V�����b�_�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�"�2�}����&����l ��h_�H���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��E���8�d�n�u�w�}�W���Y�����Rd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�d�
�&��e�}���Y���F�N�����<�n�u�u�w�}�W�������R��c1��Gڊ�&�
�l�h�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�d�1�0�E��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�E߁�
����l�N��U���u�u�u�0�3�4�L���Y���F���ʴ�
��&�g��.�(��D��ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�u�u�;�8�W���Y���F�N��U���%��
�&�w�`����-����9��Z1�N���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�=�;�:�?�/�W���Y���F�N��U���u�%��
�$�}�J���!����k>��o6��-�����n�u�w�}�Wϻ�Ӆ��V]ǻN�����'�6�&�n�]�}�W������]��D��ʥ�:�0�&�u�z�}�WϿ�&����l��^	�����u�u�'�6�$�u�������R��^	������
�!�
�$��[Ͽ�&���R��^	������
�!�d�1�0�E���Y����V��=N��U���u�3�}�}�8�u��������_	��T1�Hʴ�
�!�'�|�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9��N��U���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�g�t�^Ϫ���ƹF�N��U���%�1�;�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��X ��I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���0�4�&�2�w�/����W���F�V�����4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�N�����;�u�u�u�w�4�W�������C9��Y�����6�d�h�4��)����Y������T�����2�6�d�h�6�����
����g9��1����|�u�=�;�]�}�W���Y���R��S��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�<�(������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������R��V�����'�6�&�{�z�W�W���	����W��D�����:�u�u�'�4�.�_�������C9��P1������&�g�
�$��G�ԜY�Ʈ�T��N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�f�;���P����[��=N��U���u�u�u�%�%�<���Y����\��h�����n�u�u�u�w�8����Y���F�N�����4�,�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʴ�
�0� �;�g�a�W���&����P��h]�����
�&�<�;�1��E���	��ƹF��G1�����
�u�h�:�#���������D��R1�����
� �d�`��n�}���Y����V��Y1�I��� �
�%�'�2�)�B�������@��Y1��*��b�%�n�u�w�<�(�������Z�Y����l�6�&�
�"�l�E߁�H��ƹF�N��*���
�1�
�d�w�.����	����@�CךU���%�&�2�7�3�l�C���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z������!�9�d�d�j�<�(��������Y��D���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�f�w�.����	����@�CךU���%�&�2�7�3�l�C���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z������!�9�d�d�j�<�(��������Y��G���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�c�w�.����	����@�CךU���%�&�2�7�3�l�C���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z������!�9�d�d�j�<�(��������Y��C���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�b�w�.����	����@�CךU���%�&�2�7�3�l�C���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z������!�9�d�d�j�<�(������F��@ ��U��|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�o�}����Ӗ��P��N����u�%�&�2�5�9�F�������]9��X��U���6�&�}�%������Y����V��=N��U���u�u�u�u�w�-��������R�
N�����;�!�9�d�f�`����*����W��S�����l�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��l�W�������A	��D�X�ߊu�u�%�&�0�?���N����Z��G��U���'�6�&�}�'��(���P�����^ ךU���u�u�u�u�w�}��������lT��R��]���6�;�!�9�f�l�JϿ�&����@�
�����f�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��o�W�������A	��D�X�ߊu�u�%�&�0�?���M����Z��G��U���'�6�&�}�'��(���P�����^ ךU���u�u�u�u�w�}��������lT��R��]���6�;�!�9�f�l�JϿ�&����@�
�����l�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��n�W�������A	��D�X�ߊu�u�%�&�0�?���H����Z��G��U���'�6�&�}�'��(���P�����^ ךU���u�u�u�u�w�}��������lT��R��]���6�;�!�9�f�l�JϿ�&����@�N�����u�f�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��D���
������T��[���_�u�u�%�$�:����K�ޓ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��V��H���%�6�;�!�;�l�F������l ��_����!�u�c�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h\�U��}�%�6�;�#�1�F��DӇ��p5��D��Eʱ�"�!�u�e�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����@Ӈ��Z��G�����u�x�u�u�6���������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h]�I���4�
��3�:�m��������[��G1�����9�d�d�n�w�}����	����@��=d��U���u�%�&�2�5�9�A���
������T��[���_�u�u�%�$�:����O¹��@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9��R��]���6�;�!�9�f�l�JϿ�&����@�
�����`�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��m�����Ƽ�\��D@��X���u�4�
�<��9�(�������]9��X��U���6�&�}�%������Y����V��=N��U���u�u�u�u�w�-��������F�F��*���&�
�#�
�w�}����&����S��X����|�n�u�u�2�9��������9l�N�U���&�2�7�1�o�}����Ӗ��P��N����u�%�&�2�5�9�O߁�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������Z������!�9�d�d�j�<�(��������Y��M���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�m�6�.��������@H�d��Uʴ�
�<�
�1��e��������\������}�%��
�$�t�W�������9F�N��U���u�u�u�%�$�:����A���N��h�����#�
�u�u�'��(���Q����\��XN�\��u�u�0�1�'�2����s���F������7�1�l�d�6�.��������@H�d��Uʴ�
�<�
�1��m�(�������A	��N�����&�4�
��1�0�}���Y����]l�N��U���u�u�u�4��4�(���&����[�V�����
�#�
�u�w�-�4���
����W	��C��\��u�u�0�1�'�2����s���F������7�1�l�u�$�4�Ϯ�����F�=N��U���&�2�7�1�n���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����N�����T�����d�d�h�4������H�ƨ�D��_�\�ߊu�u�;�u�%�>���s���K�V�����&�$��
�#�m����@Ӈ��Z��G�����u�x�u�u�6�����
����g9��^�����
�&�<�;�'�2�W�������@N��h��*���
�g�|�u�w�?����Y���F��QN�����2�7�1�g�c�}����s���F�N�����<�
�&�$����������Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����9��Z1�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���
�&�$���)�E�������R��P �����&�{�x�_�w�}��������B9��h��G���8�d�
�&�>�3����Y�Ƽ�\��DF��*���
�1�
�m�]�}�W������F�N��U´�
�<�
�1��e�W������F�N��Uʴ�
�<�
�&�&��(���K����lW��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��h��*��i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�&�&��(���J����lW��V�����'�6�&�{�z�W�W���	����l��F1��*���f�3�8�d��.����	����	F��X��´�
�<�
�1��j�^���Yӄ��ZǻN��U���3�}�%�&�0�?���M�Ƹ�V�N��U���u�u�4�
�>�����*����U��D��G��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}��������V��c1��Dي�&�
�g�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�4�
�>�����*����R��D��Fʴ�&�2�u�'�4�.�Y��s���R��^	������
�!�a�1�0�F܁�
����l��TN����0�&�4�
�>�����J��ƹF��R	�����u�u�u�3��-�������� W�C��U���u�u�u�u�w�<�(���&����l5��D�*���
�f�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӇ��@��T��*���&�d�
�&��n�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<�(���&����l5��D�*���
�`�4�&�0�}����
���l�N��*���
�&�$���)�A�������R��P �����o�%�:�0�$�<�(���&����V�N�����;�u�u�u�w�4�Wǿ�&����Q�� ^�����u�u�u�u�w�}�WϿ�&����P��h=����
�&�
�`�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�d��.�(��E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϿ�&����P��h=����
�&�
�c�6�.��������@H�d��Uʴ�
�<�
�&�&��(���N����lW��V�����'�6�o�%�8�8�ǿ�&����Q��]����u�0�<�_�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y����C9��P1������&�d�
�$��A��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�F؁�
����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�d�
�$��OϿ�
����C��R��U���u�u�4�
�>�����*����_��D��M���&�2�
�'�4�g��������C9��P1����|�u�u�7�0�3�W���Y����UF��G1�����1�l�|�!�2�}�W���Y���F��G1�����0�
��&�f�����A���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�&�2�6�2��#���Hʹ��^9��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����0�
��&�f�;�������]F��X�����x�u�u�4��4�(�������@��Q��E���&�2�
�'�4�g��������C9��P1����|�u�u�7�0�3�W���Y����UF��G1�����1�f�|�!�2�}�W���Y���F��G1�����0�
��&�f�;���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�g�
�$��NϿ�
����C��R��U���u�u�4�
�>�����*����V��D��L���&�2�
�'�4�g��������C9��P1����a�_�u�u�2�4�}���Y���Z �V�����1�
�m�|�#�8�W���Y���F������6�0�
��$�o�(���&���F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�&�2�4�8�(���
����U��W��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�o�(���&����@��YN�����&�u�x�u�w�<�(���&����l5��D�*���
�e�4�&�0�����CӖ��P�������7�1�g�c�]�}�W������F�N��U´�
�<�
�1��h�^Ϫ���ƹF�N��U���%�&�2�6�2��#���K¹��^9��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���%�&�2�6�2��#���K����lW��D��ʥ�:�0�&�u�z�}�WϿ�&����P��h=�����3�8�d�4�$�:�(�������A	��D�����2�7�1�d�c�W�W�������F�N�����4�
�<�
�3��F�������9F�N��U���u�%�&�2�4�8�(���
�ԓ�@��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�'�.��������l��h��*���h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���&�2�6�0��	����������^	�����0�&�u�x�w�}��������V��c1��F���8�g�4�&�0�����CӖ��P�������7�1�d�a�]�}�W������F�N��U´�
�<�
�1��n�^Ϫ���ƹF�N��U���%�&�2�6�2��#���J����lT�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�%�$�:����&����GU��D��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C�����2�6�0�
��.�C�������@��YN�����&�u�x�u�w�<�(���&����l5��D�����f�4�&�2��/���	����@��G1�����1�g�b�_�w�}����s���F�^�����<�
�1�
�f�t����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����l ��h]��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�h����MӇ��Z��G�����u�x�u�u�6�����
����g9��1�����4�&�2�
�%�>�MϮ�������D�����l�d�_�u�w�8��ԜY���F��F��*���
�1�
�e�~�)����Y���F�N�����2�6�0�
��.�B������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�&�2�4�8�(���
�ӓ�@��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����0�
��&�a�;�������]F��X�����x�u�u�4��4�(�������@��Q��@���&�2�
�'�4�g��������C9��P1����|�u�u�7�0�3�W���Y����UF��G1�����1�c�|�!�2�}�W���Y���F��G1�����0�
��&�a�;���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�b�3�:�k�����Ƽ�\��D@��X���u�4�
�<��.����&����U��1�����
�'�6�o�'�2��������T9��S1�A�ߊu�u�0�<�]�}�W���Y���R��^	�����c�|�!�0�w�}�W���Y�����D�����
��&�b�1�0�A��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�@������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�l�3�8�o�<����Y����V��C�U���4�
�<�
�$�,�$���ʹ��^9��V�����'�6�o�%�8�8�ǿ�&����Q��^��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��M���!�0�u�u�w�}�W���YӇ��@��T��*���&�l�3�8�o�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����0�
��&�n�;���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�?����>����G9��1��*���
�g�i�u�#�-�Eځ�����l��V �����3�
�g�
�e�f�W�������`��C1�B���
�d�
�d�k�}�$���*����lW��h ��*���g�b�%�n�w�}����;����G9�� 1�����
�e�
�g�k�}��������9��h��*���d�e�%�u�8�}��������EU��^�E��|�_�u�u���$�������lW��B1�G���u�h�_�u�w�}�W���8����F��W�����f�e�"�0�w�:����&����CT�N��R��u�9�0�_�w�}�W���*����K)��h_�*؊� �g�m�%�l�}�Wϸ�&����|��X��G���
�c�
�d�k�}�$���*����lW��h ��*���g�g�%�n�w�}����;����G9��1�����;�
� �g�a�-�W������`��C1�L���2�d�d�n�w�}����;����G9��1��*��
�e�i�u�9�?����B��� ��v,��:���d�l�3�
�g��F��Y����\��h��G���d��e�n�w�}����;����G9��1�����
�c�
�g�k�}����;����G9��1�����;�
� �g�a�-�W���Y����\��h��G��e�e�e�|�]�}�W���8����F��h�����3�
�l�
�f�a�W���8����F��W��*���g�g�%�n�w�}����;����G9��Q��D݊�f�i�u�u�w�}�WϷ�&����R9��@��U²�%�3�
�f��o�G���Y�����RNךU���u�u�������N����W��G_�U���3�
��-�"���������^��G_��Hʳ�
��-� �����N����9F������d�
�
� �b�j����D���F�N��*���=�
�u�=�9�u�����ԓ�F9��1��]���h�r�r�u�;�8�}���Y���U5��C1�F���
�a�
�f�]�}�W������� 9��Q��@ފ�f�i�u�u�w�}�Wϸ�&����|��X��G���2�d�`�u�?�3�_���&����l ��[�����|�h�r�r�w�1��ԜY���F��h��D���g�3�
�a��n�}���Y����G9��1�����c�
�f�i�w�}�W���YӀ��r$��x��D���'�2�d�d�w�5��������C^��B1�D���}�|�h�r�p�}����s���F�Q=����f�`�3�
�a��D�ԜY�ƪ�l��_��@���
�c�
�f�k�}�W���Y����`9��d����b�'�2�d�d�}����Q����G��h��A���%�}�|�h�p�z�W������F�N��*���d�f�f�3��h�(��s���U5��C1�F���
�a�
�f�k�}�W���Y����]9��G��Dʢ�0�u�<�8��(�D���	����[�I�����u�u�u�u�w�;�(�������P��E��D��n�u�u�3��)�F���K����T��G]��H�ߊu�u�u�u���$�������l��h_�Eʢ�0�u�&�9�#�-�(���M�ד�N��S��D���0�&�u�u�w�}�Wϸ�&����V��B1�A���n�u�u�3��)�F���J����T��G]��H�ߊu�u�u�u���$�������l��h_�Eʢ�0�u�&�9�#�-�(���M�Г�N��S��D���0�&�u�u�w�}�Wϸ�&����V��h��@���%�n�u�u�1����I�ғ�F9��1��U��_�u�u�u�w��6���6����_��R	��F��"�0�u�&�;�)�ׁ�����l��G��U��|�0�&�u�w�}�W�������lW��hW�� ���`�%�n�u�w�;�(���H�֓�l ��]�����h�_�u�u�w�}�$���*����lW��h\�����f�g�"�0�w�.����	˹��lS��h�E���u�d�|�0�$�}�W���Y����`9��h_�*ي� �`�b�%�l�}�Wϸ�&����V��h��@���%�u�h�_�w�}�W���*����K)��h_�*؊�0�
�f�g� �8�WǷ�����lU��h�E���u�d�|�0�$�}�W���Y����`9��d����l�'�2�d�f�f�W�������lW��hY�� ���d�%�u�h�]�}�W���Y����q5��B��Cӊ�0�
�f�e� �8�Wǭ�����9��hZ�*��e�u�u�d�~�8����Y���F��d1��*��
�
� �`�b�-�L���YӀ��P��^��*���`�m�%�u�j�W�W���Y�ƪ�l'��O!��*��
�
�0�
�d�o� ���Yە��l�� 1��*���
�g�e�u�w�l�^ϻ�
��ƹF�N��&���
�g�
�
�"�h�F���B��� ��T��Gڊ�
� �`�`�'�}�J�ԜY���F��h/�����
�c�
�
�2��D��������h��F���
�b�
�g�g�}�W��PӃ��VFǻN��U����6�
�g�����A����9F������g�
� �`�c�-�W��s���F�Q=��7��� �
�c�
�2��D��������h��G���
�g�
�g�g�}�W��PӃ��VFǻN��U�������#�l�N������� S��=N��U���6�
�l�d�1��Gց�J���9F�N��U������!�f�j����H����D��F����� �f�e�%��t�J���^�Ʃ�@�N��U���3�
��-�"��Aց�&����U��d��Uʳ�
�!�l�
��(�C���	���l�N��Uʳ�
��-� ��k�(���&������YN�����8�g�3�
�e��E��Y���O��[�����u�u�u��4��N�������
9��d��Uʳ�
�!�l�
��(�C���	���l�N��Uʼ�
�9�=�
�w�5��������CQ��B1�D���}�|�h�r�p�}����s���F�Q=����
�
� �a�`�-�L���YӀ��P��1�����e�
�f�i�w�}�W���Yӏ��R
��V1����u�&�9�!�'����H����O�I�\ʰ�&�u�u�u�w�}��������9��hZ�*��_�u�u��4��N�������9��R�����u�u�u����8���H�ߓ�V��_����u�&�9�!�'����O����O�I�\ʰ�&�u�u�u�w�}�������� 9��hZ�*��_�u�u��4�����*����G��hZ��G���
�f�
�f�k�}�W���Y����V��[�����}�8�
�
�2��D��I���W����ߊu�u�u�u��%�"�������Q��1����a�n�u�u�1�����
����A��B��A؊�
� �l�d�'�}�J�ԜY���F��h��9����!�d�`�d�/���M�ƻ�V�D�����`�'�2�d�f�u�^��^���V
��d��U���u�3�
�!��.�(�������V9��h��L���%�n�u�u�1�����
����A��B��A؊�
� �l�b�'�}�J�ԜY���F��P1�Lʢ�0�u�&�9�#�-�@�������
N��S��D���0�&�u�u�w�}�Wϸ�&����R��d�����0�a�
�
�"�d�F���B��� ��T������'�6� �2�i�(ց�����l��S��U���u�u�'�2�f�d� ���Yە��l��W�����a�c�e�u�w�l�^ϻ�
��ƹF�N��&���
�4�0��%�>����M����U��Y��F�ߊu�u��6��<��������A��1��*���
�f�i�u�w�}�W�������S��_��]���6�;�d�d��8�(��L���F�G�����_�u�u�u�w���������G��C��*���g�3�
�f��n�}���Y����G9��D�����!�'�
�l�f�;�(��&���FǻN��U����-� ��9�(�(��&����T9��]�����}�'�6�;�f�l�(���&����V�
N��R���9�0�_�u�w�}�W�������@��C�����
�l�3�
�c��D�ԜY�ƪ�l��t��*��� �!�'�
�n�o����A˹��Z�=N��U���u�0�
�`�w�5��������CW��E��D��}�|�h�r�p�}����s���F�Q=�����&�
�!� �#�/�(���H����
^��G]�U���3�
�!��$���������_��h��L���%�u�h�_�w�}�W�������F��R �����!�%�b�'�0�l�F���P���A�R��U���u�u�u�3��)�4���&����P��R1�*؊� �l�m�%�l�}�Wϸ�&����R��d�����0�a�
�
�"�l�G݁�J���9F�N��U���-� ��;�"��@ځ�&����R�������0�
�8�d��8�(��O���F�G�����_�u�u�u�w���������G��C��*���f�3�
�l��n�}���Y����G9��D�����!�'�
�l�1��Cށ�J���9F�N��U���
�`�u�=�9�u����&����U��^��H��r�u�9�0�]�}�W���Y����P��=N��U���6�
�4�0��/��������9��h_�L���u�h�_�u�w�}�W���&����D��F��*���1�
�a�'�0�l�G���P���A�R��U���u�u�u�3��)�4���&����P��R1�*���l�m�%�n�w�}��������V9��E�� ���`�
�
� �f�l�(��E��ƹF�N�����c�u�=�;��8�(���Hƹ��T9��\��\��r�r�u�9�2�W�W���Y�ƪ�l��t��*��� �!�'�
�a�l����I�ߓ� ]ǻN��&���
�4�0��%�>����LŹ��U��\�����h�_�u�u�w�}�$���,����|��Y��F���2�d�a�u�?�3�_���&����9��P1�D���|�h�r�r�w�1��ԜY���F��h��6���
�!� �!�%��A�������P��UךU����6�
�4�2���������9��Q��E���%�u�h�_�w�}�W�������F��R �����!�%�l�'�0�l�E���P���A�R��U���u�u�u�3��)�4���&����P��R1�*ي� �d�g�
�d�W�W���*����p��h=�� ���'�
�c�3��i�(��E��ƹF�N��&��� ��;� ��j�(܁�����U��_��]���
�
�0�
�d�n�G���Y�����RNךU���u�u�0�
�b�f�W�������A��~ �����
�;�
�:�%�8�A�������S��N�U���u�u�u�4��2�����ԓ���YN����� �d�a�%��t�J���^�Ʃ�@�N��U���3�
�!��$���������P��h��*��c�_�u�u��)����0����]��V ��6���6�
�
� �f�i�(��E��ƹF�N�����;�!�9�f��}����Q����U��W��G��u�u�d�|�2�.�W���Y��� ��T������'�6� �2�i�(ց�����V��N�����0�8�
�;��3��������A�� 1��*��f�%�u�h�]�}�W���Y����\��h��G��"�0�u�2�'�;�(��&���F�_��U���0�_�u�u�w�}�$���&����l5��B�����g�l�'�2�f�h�L���YӀ��K'��N!��*���
�l�
� �`�h����DӔ��lW��d��Uʳ�
���g��)�F���J����
T��G]��H�ߊu�u�u�u��%�"�������Q��Q��Eߊ�d�"�0�u�$�1����J����
T��G\��\��r�r�u�9�2�W�W���Y�ƾ�T9��UךU����-� ��9�(�(��&����S��N�U���0� �!�d��(�O���	��ƹF��d1�� ���;� �
�b��3����/�ד�F9��1��U��&�1�9�2�4�+����Q����T�������!�&�3�
�e��D���Y����T�������!�9�f�
���1���P��ƹF��d1�� ���;� �
�b��3����	����l^��h�I���u�u�u�u�%�)�E�������G9��D�� ��l�%�u�=�9�u��������U��_��G��u�u�d�|�2�.�W���Y�����h��A���
�l�
�f�]�}�W��Y����U��]��ʴ�&�2�u�'�4�.�Y��s���T��Q��Eي�0�4�&�2��/���	����@��G1��Yʴ�
�<�
�&�&��(���&����J��G1�����0�
��&�c�;���Y����Z��D��&���!�
�&�
�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t��������]��[����h�4�
�<��.����&����U��G�����%�6�;�!�;�:���DӇ��@��T��*���&�`�3�8�c�t�^Ϫ���ƹF�N��U���'�
� �d�d�>�W������]��[����_�u�u�u�w�1��ԜY���F�N�����
�e�
�0�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R�����u�2�%�3��m�(��E�ƪ�l��_��A���2�d�l�n�w�}�������� 9��R�����!�d�e�a�%�:�F��B���F�	��*���d�a�:�6�3�}����Ӗ��P��N����u�'�
� �f�i��������@��h����%�:�0�&�6�����
����g9��1����u�%�&�2�4�8�(���
�Փ�@��N��*���
�&�$���)�G���������h��D���1�8�'�4��8�(��K�ƭ�l��h�����
�!�d�3�:�o�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1�����0�
��&�e�����I�ƭ�WF��R����d�1�8�'�6�����M�����T�����d�e�|�u�?�3�}���Y���F�P�����d�
�%�:�2�a�W�������l
��hZ�U���u�u�0�&�1�u�_�������l
��^��U���%�&�2�6�2��#���J����lT�X�����:�&�
�:�>��W���	����l��F1��*���e�3�8�d�~�t����Y���F�N��U���
� �d�a�8�>����DӇ��P	��C1��@��_�u�u�u�w�1����Q����\��h�����u�u�%�&�0�>����-����l ��h_��U���;�_�u�u�w�}�W�������lW��h�����i�u�%�6�9�)����K���F�N�����u�u�u�u�w�}��������9��T��U��w���w�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�ƫ�C9��h_�*��4�&�2�u�%�>���T���F��G1��*��
�e�4�&�0�����CӖ��P�������4�d�u�%�$�:����&����GT��D��Yʴ�
�<�
�&�&��(���&����J��d1��*���0��'�6�"�8�C݁�&����R��B��&���
�4�0��%�>����M����A��Z�Yʴ�
�<�
�&�&��(���I����lW�������6�0�
��$�o�(���&���F�U�����u�u�u�<�w�u��������\��h_��U���&�2�6�0��	���&����V����ߊu�u�u�u�w�}��������l��S��&���
�4�0��%�>����M����A��Z�N���u�u�u�0�$�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����֓�@��G�����u�u�u�u�w�}�WϹ�	����W��G^��Hʳ�
�!��&��)��������l_��B1�A���n�u�u�u�w�8����Q�έ�l��D�����
�u�u�%�$�:����&����GT��D��\ʺ�u�4�
�:�$�����&���R��^	������
�!�
�$��^�������9F�N��U���u�'�
� �f�i����Dӏ��R
��V1����u�u�u�9�2�W�W���Y���F��G1��*��
�e�i�u���/���!����k>��o6��-�������l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����A��B1�A���u�&�<�;�'�2����Y��ƹF��E�� ��a�%�
�&�>�3����Y�Ƽ�\��DF��*���
�&�$���)�(���&����C9��P1������&�f�3�:�o�W���
����@��d:�����3�8�d�y�6�����
����g9��_�����e�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`��������V��c1��Gڊ�&�
�l�|�#�8�W���Y���F�	��*���d�a�%�u�j�<�(���
���� T��qV�E��_�u�u�u�w�1����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���}�%�6�;�#�1����H����C9��P1������&�f�3�:�o�W���Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���!�0�u�u�w�}�W���YӁ��l ��_�����h�4�
�:�$�����I���F�N�����u�u�u�u�w�}��������9��R��W���������/���!����k>��o6��W�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�/�(���H�֓�C��RN�����u�'�6�&�y�p�}���Y����U��^�����0�4�&�2��/���	����@��G1�����0�
��&�e�;���Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�*���
�l�u�0��0�E�������T��E��D��y�4�
�<��.����&����l ��h\����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�4�1�}�2����H����\��Y1����l�u�u�%�4�3����H���F��R ��U���u�u�u�u�0�-����Kù��P	��R�����:�&�
�#��f�W���Y����_��F�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�8�}��������_	��T1�Hʴ�
�<�
�&�&��(���I����lW��G�����_�u�u�u�w�}�W���&����V��G����u�%�6�;�#�1�B��s���F�R�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�W������F�N��Uʲ�%�3�
�g��-����E�ƭ�l��D��ߊ�n�u�u�u�w�8����Y���F�N����� �d�e�:�4�9�W��[����kD��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�2�%�3��o�(������]F��X�����x�u�u�2�'�;�(��&�֓�@��Y1�����u�'�6�&���6���6����_��R	��F��u�%�&�2�4�8�(���
�ԓ�@��N��*���
�&�$���)�(���&����C9��P1������&�g�
�$��N���*����p��h=�� ���'�
�l�l�1��G���	����`9��h-�����'�6� �0�c��(���&����F��h��*���$��
�!�f�;���P�����^ ךU���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�F�������F��R ��U���u�u�u�u�0�-����Kù��Z�Q=�����&�
�!� �#�/�(���@����lW��UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	���&����_����ߊu�u�u�u�w�}��������l��S��&���
�4�0��%�>����Mʹ��U��^����u�u�u�u�2�.����Q����\��h�����u�u�%�&�0�>����-����l ��h_�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�^Ϫ���ƹF�N��U���'�
� �d�g�-�W������`��C1�L���2�d�d�n�w�}�W�������9F�N��U���u�'�
� �f�m����D�Ĕ�k>��o6��-���������/���!����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʲ�%�3�
�g��l�����Ƽ�\��D@��X���u�2�%�3��o�(�������]9��X��U���6�&�}�%�$�:����&����GT��D��Yʴ�
�<�
�&�&��(���&����J��G1�����0�
��&�e�����@�ƭ�l��h�����
�!�d�3�:�o�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��h��*���$��
�!�g�;���P�Ƹ�V�N��U���u�u�2�%�1��E߁�H���R��X ��*���g�f�m�e�g�f�W���Y����_��F�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�8�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��EN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�e�~�}����s���F�N�����3�
�g�
�f�a�W�������l
��1����u�u�u�9�2�W�W���Y���F��G1��*��
�d�i�u���/���!����k>��o6��-�������l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����A��B1�@���6�1�u�&�>�3�������KǻN����� �d�`�:�4�9�(�������A	��N�����&�4�
�<��.����&����U��B�����2�6�0�
��.�E߁�
����F��[1����
�0�:�2�9�/���H����C9��P1������&�g�
�$��G�ԜY�Ʈ�T��N��U���<�u�}�4��2��������F�V�����&�$��
�#�l����K����]�D�����d�
�0�:�0�3����H����F��h�����#�
�|�|�#�8�W���Y���F�	��*���d�`�:�6�3�}�JϿ�&����G9��1����u�u�u�9�>�}�_ǿ�&����G9��P��D��4�
�<�
�$�,�$�������^9����]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�n�t�W������F�N��Uʲ�%�3�
�g��-����E�ƭ�l��D��ߊ�n�u�u�u�w�8����Y���F�N����� �d�`�:�4�9�W��[����kD��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�2�%�3��o�(������]F��X�����x�u�u�2�'�;�(��&�֓�@��Y1�����u�'�6�&��-��������`2��C\�����y�4�
�<��.����&����l ��h_�U���6�
�4�0��/��������9��h_�L���y�3�
�!��.�(�������V9��hV�����a�c�u�%�$�:����&����GT��Q��G���3�
��-�"��(���K�ѓ� OǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����ד�@��G�����u�u�u�u�w�}�WϹ�	����T��G^��Hʳ�
�!��&��)��������l^��R	��A��_�u�u�u�w�1����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y����U��[��E��u��6�
�6�8�$�������lS��1��*��l�%�n�u�w�}�Wϻ�
�����T�����2�6�d�h�6�����
����g9��1����|�!�0�u�w�}�W���Y����A��B1�@���u�h�3�
��%����&����Q��UךU���u�u�9�0�]�}�W���Y���T��Q��Gߊ�e�i�u����/���!����k>��o6��-������n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӁ��l ��\�����&�<�;�%�8�8����T�����h��D���%�
�&�<�9�-����Y����V��V�����&�$��
�#�����UӇ��@��T��*���&�g�
�&��d�W���
����@��d:�����3�8�g�y�1��5�������
9��Q��B؊�f�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`��������V��c1��Gۊ�&�
�e�|�#�8�W���Y���F�	��*���d�`�%�u�j�<�(���
���� T��d��U���u�0�&�3��<�(���
����T��N�����<�
�&�$����������
O�C��U���u�u�u�u�w�:����&����CW�
N��*���&�
�#�g�d�e�G��B���F������}�%�6�;�#�1����H����C9��P1������&�g�3�:�l�^Ϫ���ƹF�N��U���'�
� �d�b�-�W������`��C1�L���3�
�b�
�d�W�W���Y�Ʃ�@�N��U���u�u�2�%�1��Eځ�H���>��o6��-���������/���!����]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�'�
� �f�i����
������T��[���_�u�u�'��(�F���	ù��@��h����%�:�0�&�6�����
����g9��1����u�8�
�
�"�o�G���UӒ��lT��R	��F��u�%�&�2�4�8�(���
�Փ�@��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����l ��h\��U���;�_�u�u�w�}�W�������lW��h�I���8�
�
�0��n�C�ԜY���F��D��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}����s���F�N�����3�
�f�
�g�a�W���&����lT��h����u�u�u�9�2�W�W���Y���F��G1��*��
�e�i�u��f�W���Y����]��QU��U���0�1�%�:�2�.�}���YӁ��l ��]�����h�}�'�
�"�l�C���Y����T��Q��Dފ�g�n�_�u�w�p��������
9�������%�:�0�&�w�p�W�������F9��1��*���<�;�%�:�w�}����
�έ�l��h�����
�!�
�&��q����Hǹ��lT��h�U���
�a�'�2�f�i�[Ͽ�&����P��h=�����3�8�g�_�w�}����s���F�^��]���6�;�!�9�0�>�F������T9��R��!���f�3�8�g�~�)����Y���F�N����� �d�l�%�w�`����Hǹ��T9��Y�U���u�u�0�&�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O�C��U���u�u�u�u�w�:����&����CV�
N����
� �g�`�'�f�W���Y����_��=N��U���u�u�u�'��(�F���	���D��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���2�%�3�
�d��E��Yہ��l ��]�����;�u�'�
�"�l�G���P��ƹF�N�����
�a�
�e�6�.��������@H�d��Uʲ�%�3�
�a��m��������\������}�%�&�2�4�8�(���
����U��W����f�
� �d�o��E�������l��h_�B���%�&�2�6�2��#���K¹��^9��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y����U��Z��E��u�8�
�f�%�:�F��B���F������}�%�6�;�#�1����H����C9��P1������&�g�
�$��N�������9F�N��U���u�'�
� �f�i����DӒ��lU��Q��E���%�n�u�u�w�}����Y���F�N��U���
� �d�a�'�}�J���[���F�N��ʼ�n�_�u�u�9�}����
��ƓF�P�����a�
�g�i�w�:����&����CV��Y
����� �d�a�%�~�W�W���T�ƫ�C9��h_�*��4�&�2�u�%�>���T���F��G1��*��
�e�4�&�0�����CӖ��P�������6�0�
��$�o�(���&���G��V�� ��a�
�g�u�:��O�������J��G1�����0�
��&�e�����I���F��P��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�Eށ�
����O��_�����u�u�u�u�w�/�(���H�ߓ�F���*���'�2�d�l�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��Gڊ�&�
�l�|�#�8�W���Y���F�	��*���d�l�%�u�j�)���&����R��G\�U���u�u�0�&�w�}�W���Y�����h��D���%�u�h�w�u�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����U��W��G��u�2�%�3��i�(������A��B1�E���|�_�u�u�z�}��������l��V�����'�6�&�{�z�W�W�������lW��h�����2�
�'�6�m�-����
ۇ��@��T��*���&�g�
�&��d�W���&�Փ�F9��Y��G���8�
�f�'�0�l�G������T9��R��!���g�
�&�
�g�W�W�������F�N�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��G�������9F�N��U���u�'�
� �f�i����DӒ��lR��E��D��n�u�u�u�w�8����Qۇ��P	��C1�����d�h�4�
�>�����*����V��D��L���!�0�u�u�w�}�W���YӁ��l ��[�����h�!�%�a��(�F��&����F�N�����u�u�u�u�w�}�WϹ�	����S��G^��H���w�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�/�(���H�ғ�F�F�����
�`�
�e�6�9��������9��UװU���x�u�'�
�"�d�(�������]F��X�����x�u�u�2�'�;�(�������@��h����%�:�0�&�6�����
����g9��1����u�%�6�y�6�����
����g9��1����u�%�&�2�4�8�(���
�Փ�@��N��*���
�&�$���)�D���������D�����
��&�g��.�(��Y����Z��D��&���!�d�3�8�e�t�W�������9F�N��U���}�}�%�6�9�)���������D�����
��&�d�1�0�G���ӈ��N��h�����:�<�
�u�w�-����Y���R��X ��*���<�
�u�u�'�.��������l��h��*���:�u�4�
�8�.�(�������F��h��*���$��
�!��.�(�������C9��Y�����6�d�h�4��4�(�������@��h��*��u�'�}�%�4�3��������[��G1�����0�
��&�e�����@�ƣ�N��h�����:�<�
�u�w�-��������`2��C\�����g�|�|�!�2�}�W���Y���F��E�� ��
�0�i�u�'�>��������lV��N��U���0�&�u�u�w�}�W���YӁ��l ��W����u�%�6�;�#�1����H���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����3�
�l�:�4�9�W�������A	��D�X�ߊu�u�'�
�"�d�(�������@��Y1�����u�'�6�&��-��������`2��CY�����y�4�
�<��.����&����U��B�����2�6�0�
��.�F߁�
������D�����
��&�d��.�(��Y����Z��D��&���!�b�3�8�f�t�W�������9F�N��U���}�}�%�6�9�)���������D�����
��&�d��.�(��Y���R��X ��*���<�
�u�u�'�.��������l�� 1����|�|�!�0�w�}�W���Y�����h��Lӊ�%�:�0�i�w�-��������lW��N��U���0�&�3�}��-��������Z��S�����2�6�0�
��.�@������\�V�����
�:�<�
�w�}��������B9��h��*���
�|�:�u�6�����&����P9��
N��*���
�&�$���)�G������F��R ��U���u�u�u�u�0�-����@����\��S�����;�!�9�g�g�W�W���Y�Ʃ�@�N��U���u�u�2�%�1��N�������[�o6�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�%����&����@��YN�����&�u�x�u�w�:����&�ߓ�9��D��*���6�o�%�:�2�.����H���A��X�U���6�
�l�a�%�:�F��UӇ��@��T��*���&�b�3�8�a�}�$���,����|��Y��F���2�d�a�y�6�����
����g9��1����u�%�&�2�4�8�(���
����U��B�����2�6�0�
��.�Fہ�
����F��h��*���$��
�!�`�;���P�����^ ךU���u�u�3�}�6�����&����P9��
N��*���
�&�$���)�C�������F��R ��U���u�u�u�u�0�-����@����[��d1�� ���;� �
�b������M����F�N�����3�}�4�
�8�.�(�������F��h��*���$��
�!�g�;���PӒ��]FǻN��U���u�u�'�
�"�d�(��E�ƾ�T9��UךU���u�u�9�<�w�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��EN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�c�~�}����s���F�N�����3�
�l�%�w�`����H����F�N�����3�}�4�
�8�.�(�������F��h��*���$��
�!��.�(���Y����l�N��U���u�2�%�3��d����DӀ��P��1�����d�m�n�u�w�}�Wϻ�
��ƹF�N��U���'�
� �l��m�K���!����k>��o6��-���������/���B���F���U���u�u�u�0�3�-����
��ƓF�C����� �l�
�d�6�.��������@H�d��Uʲ�%�3�
�l�'���������PF��G�����<�
�4�
�{�/���@�ƪ�l��\��@���2�d�m�y�1��6���6����W��R	��A��u�%�&�2�4�8�(���
�ѓ�@��N��*���
�&�$���)�(���&����C9��P1������&�d�
�$��[Ͽ�&����P��h=����
�&�
�f�w�-��������`2��C_�����d�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�5��ԜY���F�N�����
�l�%�u�j�/���@���F�N�����}�}�%�6�9�)���������D�����
��&�d��.�(�������C9��Y�����6�d�h�4��4�(�������@��h��*��|�u�=�;�]�}�W���Y���T��Q��L���u�h�3�
���8���H�ד�V��]����u�u�u�9�>�}�_�������l
��^��U���%�&�2�6�2��#���N����lP����ߊu�u�u�u�w�}��������CW�
N��*���
�n�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��Q��F���!�0�u�u�w�}�W���YӁ��l ��W��D��u��6�
�e��(���&����l�N��Uʰ�&�u�u�u�w�}�W�������F9��h�I���������/���!����k>��o6��-���n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�>�0�@���&����CT�
N��Wʢ�0�u�!�%�d����N����F��h�����#�
�|�0�$�}�F��Y����P��h ��*���c�g�%�u�j�u����&����R��N��ʴ�
�:�&�
�!��^�ԜY�ƥ�^��B1�E���u�h�w�w� �8�WǪ�	����U�� ]��F��4�
�:�&��+�(�������V�=N��U���%�;�!�3��i�(��E����P��Q��Mڊ�g�-�'�4��2����¹��l�N��*���=�
�
�:�>�)����Nù��Z�^ �����
�n�u�u�;�>�!�������
9��R��������!��9�F�������9��\�X��1�"�!�u�~�W�W�������9��h_�D���u�h�%��;��(���H����CW�N�����u�f�n�u�w�1����J����V��h�I���
�4�g�d�1��G���	����K�
�����e�n�u�u�;�>�!�������T��N�U���4�g�g�3��m�O���Q����\��XN�\�ߊu�u�:�
�����H����Z�G1��؊�
� �d�l��l�E���Y�ƨ�D��^����u�:�
�
��(�F��&���F��a��*ي� �d�`�
�f�n�W������ O��N������b�3�
�f�n����DӖ��R
��1��*��l�%�}�f�z�l��������l�N�����3�
�a�
�c�a�W�������|��v
��D���3�
�a�
�f�n�W������ O��N�����0�d�3�
�d��D��Y���F������!�9�f�`� �8�WǷ�����lU��h�E���u�d�|�0�$�}�W���Y����C9��Y�����a�_�u�u�2����&����l ��\�*��i�u�!�
�8�4�(�������V��RF�����0�}� �
�2�)���&����V9��D��*���
�a�e�y�~�f�W�������_T��B1�@���u�h�_�u�w�}�W���*����R��T��*���c�l�%�u�?�3�_�������U��Y��G��u�u�d�|�2�.�W���Y�����d�����g�
�f�_�w�}��������G9��D�� ��l�%�u�h�]�}�W���Y����\��h��*���=�;�}�0��0�O���&����CT�N��R��u�9�0�_�w�}�W���	����@��A]��N���u�;�"�0��(�A���	���l�N��Uʴ�
�:�&�
�!��W����ο�_9��GY�� ��d�%�}�|�j�z�P������F�N�����:�&�
�#��f�W�������@W��B1�Lߊ�g�i�u�e�w�5��������9��h_�F���u�u�%�6�9�)����?����_��_�����u�:�9�&��(�E���	���D�������8�
�e�3��o�(��DӇ��P	��C1��M���|�0�&�u�f�f�W�������@R��B1�C���u�h�w�w� �8�WǪ�	����U��Z��A��4�
�:�&��+�(���Y����D��d��Uʻ�!�=�`�3��n�(��E���F��R �����g�
� �f�e�-�W���	����@��AV��3���9�0�w�w�]�}�W�������U��Y�����h�w�w�"�2�}����/�ԓ�F9��_��A��4�
�:�&��+�(���Y����D��d��Uʻ�!�=�m�3��l�C���Y���D��_��]���
�
�
� �f�m�(��DӇ��P	��C1��M���|�0�&�u�f�f�W�������@9��h_�*��i�u�e�u�?�3�_���&����R��N�����:�&�
�#���W�������l�N�����d�3�
�g�f�-�W��[����[����*���
� �d�b��l�JϿ�&����G9��]��\ʰ�&�u�e�n�w�}�����ԓ�F9��1��U��w�w�"�0�w�)���&���� _��N�����:�&�
�#�d�m�W�������l�N�����a�3�
�g��o�K���H�ƻ�V�C��Gڊ� �g�a�%�w�}��������ET��G�����w�w�_�u�w�2����&����V��N�U��u�=�;�}�:��E���&����CW������!�9�g�
�~�8����I��ƹF��X��܊� �d�b�
�e�a�W��Y����N��T1��F���
�e�d�%�w�}��������ET��G�����w�w�_�u�w�2����&����R��G\��H���w�"�0�u�;�>�!�������T��N�����:�&�
�#�d�m�W�������l�N�����
� �d�a�'�}�J���[ӑ��]F��Z��*���d�a�%�u�w�-�������� 9�������w�_�u�u�%�>����Hǹ��lP��h�I���<�8�b�3��j�(������V��B1�C���|�_�u�u�%�>��������9��R��]���
�8�b�3��h�(���ƿ�_9��G\�� ��d�%�|�_�w�}�����ԓ�F9��1��U��}�'�6�;��(�A���	�ƣ�	��T��D���
�f�
�g�l�}�Wϱ�&����l ��_�����h�}�0�
�:�e����I¹��	��D�����
� �a�c�'�t�}���Y����`��X��F���<�0�4�&�0����@����[�N��U���;�"�0�g�1��Cځ�Jӑ��]F��E1�����3�
�`�
�e�m�W���H����_��=N��U���u�0��9��(�A���	��ƹF��B�����0�!�f�"�>�8��������lW��1��U��_�u�u�u�w�8�(���K����lW��1��U���;�}�0�
�:�o�F�������]9��P1�D���|�h�r�r�w�1��ԜY���F��h��ۊ�;��;�0�6�9�4�������9��h_�@���n�u�u�:�#���������D��R1�����
� �d�`��n�K���Y���F��R����
� �d�`��n� ���Yە��l��^�����'�4�
�0��i�@��Y���O��[�����u�u�u��#�/�F���&����V9��S1�����
�
� �d�c��D�ԜY�ƣ�G9��R�����
�'�!�
�$�4����&����l��S��U���u�u�&�9�#�-�G���&����l��@��U¦�9�!�%�l��8��������lW��F�U���d�|�0�&�w�}�W���YӀ��G��1��*���2�
�;�
�8�/��������U��UךU���
�d�b�d�1��B؁�J���9F�N��U���6�;�!�9�e��W����θ�C9��h��M���%�}�|�h�p�z�W������F�N�����d�3�
�`��l�}���Y����@��h_�����l�
�`�i�w�;�(���=����l'��h_�*���b�`�%�}�f�9� ���Y���F��G1�*���m�`�%�|�]�}�W�������l��B1�@���u�h�}�%�4�3����KŹ��F��T1�����a�
�a�n�w�}��������U��]�����h�3�
�!��.�(�������V9��hW�� ��a�%�n�u�w�-�!���&����lW��1��U��3�
�!��$���������_��h��D��
�f�_�u�w�����J����W��h�I����6�
�4�2���������9��Q��E���%�n�u�u�%�)�E�������G9��D�� ��l�%�u�h�]�}�W���Y����\��h��@���e�"�0�u�#�-����H����lQ��h�E���u�d�|�0�$�}�W���Y����C9��Y����
�e�n�u�w�/��������Q��G]��H�ߊu�u�u�u�'�>��������V�������8�
�
�
�d�;�(��&���F�_��U���0�_�u�u�w�}��������EW��Z�N���u�'�#�3��e�(��E����\	��O)��:���d�a�'�2�f�k�W���Y����\��h��*���_�u�u�0��0�F߁�����l��S�����b�
�
�
�"�j�D���Y����@��C��*���m�`�%�|�]�}�W���&����9��hW�*��i�u�d�u�?�3�_���������C1�@���
�%�,�0�1��F؁�J����C9��Y����
�a�e�u�;�8�U���s���@��C��G���
�d�
�g�k�}�F������U5��z;��G���!�d�`�<��-��������9��S�����;�!�9�d��m�^ϻ�
���]ǻN�����8�d�
�0�8�:����&����CT�
N�����8�c�1�8�%�<�(���M�ғ�F����*Ҋ� �f�d�%�~�W�W�������CW��Q��Gۊ�g�i�u�&�;�)��������
9�������!�%�g�3��l�(��B�����h��D���1�8�'�4��(�@���	���N��h��ۊ�a�3�
�m��o��������l ��V�����_�u�u�0��0�F�������T��Q��G݊�g�i�u�&�;�)���&����A��h��B���%�u�'�!�'�e����@¹��]ǻN�����8�d�
� �a�e����D�ή�\
��p+�� ���c�
�0�
�d�n��������]	��Q��L؊�g�n�u�u�$�1����L����V��G\��H���8�
�g�3��e�(������V
��Z�*���c�m�%�|�]�}�W���&����9��hY�*��i�u�&�9�#�-�Cށ�����R��B1�L���u�:�u�%�4�3����H���9F���*���d�
� �b�f�-�W��Q����9��h]�*��4�1�&�9�#�-�A���&����CT�=N��U���
�8�d�
�"�j�D���Y���@��C��AҊ�0�:�2�;�1��E؁�KӞ����T�����d�d�n�u�w�.����	����W��E	��*���d�l�
�g�k�}��������9�������d�
�0�:�0�3����I�ѓ�O��N�����!�%�l�3��n�(��E����^��h��F���%�u�;�u�2����&���� U��G�U���&�9�!�%��(�C���	���N��Z�� ��e�%�u�:�w�-��������lW�=N��U���
�8�g�d�3�0����&����S��G\��H���'�
� �d�n�-�W�������9��Z����� �d�g�
�e�f�W���
����^��h��D��
�f�i�u�w�}�W�������]��[�*ݓ�e�e�e�"�2�}����HĹ��^	��V �����a�g�e�u�w�l�^ϻ�
��ƹF�N�����;�!�9�f���G��I���F��[1����
�0�:�2�9�;�(��M����[�P�����`�
�g�:�w�0�(�������T��Q��D���%�|�_�u�w�8�(���K¹��lW��1��U��_�u�u�u�w�-��������9��t^�E���=�;�}�8��h��������A��Z�]���h�r�r�u�;�8�}���Y���R��X ��*���g�f�m�e�g�f�W���
����^��h
�����;�3�
�m��o�K���
����^��h
�����;�3�
�c��o��������U��Y��G��u�u�&�9�#�-�E���&����l��S��U���u�u�4�
�8�.�(���K�ъ�V��N�����!�%�f�
�2�2��������V��G��U��|�0�&�u�w�}�W�������]��[�*ٓ�e�e�e�_�w�}�����ԓ�F9��1��U��}�0�
� �d�k�����ƿ�_9��G_�� ��`�%�|�_�w�}�����Փ�F9��1��U��}�8�
�
�"�n�@���Y����@��C�����b�
�g�n�w�}��������U��Y��F��u�u�u�u�w�/��������Q��G]�����}�8�
�
��(�@���	����[�I�����u�u�u�u�w�<�(���
����S��^�U���&�9�!�%��(�C���	���N��[1�����1�8�'�4��(�C���	�ƴ�AF��h�����#�
�|�_�w�}�����Г�V��P�����f�
�g�i�w�4��������l��X����� �f�c�%�~�W�W�������CP��B1�C���u�h�}�:�;�%�2�������l��h_�Fʴ�1�<�8�
�8����I����l�N�����%�
� �a�f�-�W��Q����9��h]�*��4�1�&�9�#�-�(���M�Г�O��N�����!�%�
� �b�l����D�θ�C9��Q��Eي�g�4�1�&�;�)�ځ�����l��d��Uʦ�9�!�%�
�"�e�B���Y���G��^1�����c�
�g�-�%�<�(���
����9��d��Uʦ�9�!�%�3��j�(��E����V
��Z�*���:�2�;�3��k�(������C9��Y�����d�n�u�u�#�-�F߁�����l��S��&�����!�d�n�o��������lT��h�F���:�;�:�g�~�W�W�������l ��X�����h�}�7�:������&����A��]�U���'�
� �d�n�-�^�������F9��1��\�ߊu�u�8�
�e�;�(��&���F�N�����!�%�d�
�"�n�C���Y�ƭ�l��D��ي�|�0�&�u�g�f�W������� 9��h\�*��i�u�������@�ԓ�\9��C1��*��
�d�g�u�w�}�������9F���*���3�
�`�
�e�a�Wǰ�����l ��Z�����'�;�!�=�e�;�(��&���9F���*���1�8�'�4��(�F��&���F��Z��*���3�
�e�`�'�}��������ZW��1��*��d�%�|�_�w�}����N����^��G]��H���8�
�d�3��j�(��_Ӗ��S��1��*���
�f�n�u�w�)���&����R��N�U������!�#���������l��^�����:�g�|�_�w�}����&����R��N�U���4�%�4�d�#���������l��]��U���:�;�:�e�l�}�WϪ�	����U��Z��D��u�����)��������lT��h�G���u�u�:�;�8�m�L���YӒ��lT��Q��E؊�a�i�u����8���K����Z��Q��LҊ�d�f�u�:�9�2�E���s���G��\�� ��g�%�u�h�1��5�������G	��Y�� ��m�%�}�f�z�l��������l�N����
� �f�m�'�}�J�������9��h]�*��:�u�:�9�$����O����l�N����
� �f�c�'�}�J�������9��h]�*��:�u�:�9�$����M����l�N����
�0�:�2�9�;�(��A����[�C�����
� �d�d��o��������l��X�� ��g�
�g�n�w�}����Kƹ��lU��h�I���!�%�g�
�"�n�O���Y����G��Z�� ��c�%�|�_�w�}����N���� Q��G]��H���:�9�-���)�F������� P��N�����
�f�
�g�l�}�WϪ�	����U��_��G��u�!�%�f�1��Dց�KӉ��G��1��*��
�g�n�u�w�)���&����S��N�U���u�u�u�4��2����˹����YN�����
� �m�l�'�u�^��^���V
��d��U���u�4�
�:�$��ׁ�B�����h\�� ��e�%�u�h��2��������9�������=�
� �d�o�-�^�ԜY�Ƹ�C9��h��M���%�u�h�3���;���6����S��Y1�����d�3�
�f��o�O��Hӂ��]��G�U���!�%�f�
�"�e�@���Y���F�N�����g�
� �m�b�-�W����θ�C9��h��M���%�}�|�h�p�z�W������F�N����
� �m�f�'�f�W�������9��hX�*��i�u�7�:������&����A��]�U���'�
� �d�n�-�^�ԜY�Ƹ�C9��h
�����;�3�
�d�n�-�W��Q����Z9��h��D��
�g�4�1�#�-����&�ѓ�F9��]��G��u�u�!�%�d����Aƹ��Z� �����
� �d�b��o��������9��h_�F���|�_�u�u�:��O���&����l��S�����=�m�3�
�f�m����ӈ��_��h��D��
�g�n�u�w�)��������
9��R��W���"�0�u�&�0�8�_���������C1�@���
�-�
�
��(�O���	�����Y�����:�&�
�#�c��^������D��N�����a�
� �d�g��E��Yۈ��A��h��D��
�g�:�u�8�1�ށ�����9��UךU���8�
�
� �o�h����D������YN�����1�3�
���o�8���H�ӓ�]9��G1��D���
�f�
�g�w�}����ۇ��P	��C1��Fފ�|�u�9�0�u��}���Y����_��h�� ��f�%�u�h�u�� ���Yۊ��l0��B1�L���u�u�%�6�9�)����?����_��^�����u�8�
�
�"�n�F���Y���D��_��]���
�d�3�
�a��C������]��[��@���9�0�w�w�]�}�W���&ʹ��lU��h�I���d�u�=�;��0�(�������9��S�����;�!�9�f�a�}����[����F�C�����b�
�a�i�w�3�����ד�\9��C1��*��
�d�f�u�8�3���P���F��G1��ۊ�`�3�
�e�f�-�W��[����[����*���
� �d�`��l�JϿ�&����G9��]��\ʰ�&�u�d�n�w�}��������U��[�����h�w�w�"�2�}����/�ԓ�F9��_��A��4�
�:�&��+�(���Y����D��d��Uʡ�%�<�<�
�a�;�(��K����[�L�����}�:�
�
��(�F��&�����T�����g�
�|�0�$�}�F��Y����^��h�����d�c�%�u�j��Uϩ�����\��hZ�� ��e�
�a�h�6�����&����u �R��U��n�u�u�!�'�4�؁�N����W��h�I���e�u�=�;��2�(���&����Q��G_��U���6�;�!�9�e��^ϻ�
���]ǻN�����
�b�3�
�f�j����D������YN�����
�
� �d�a��C������]��[��3���0�&�u�e�l�}�WϪ�	����lW��Q��Cӊ�g�i�u�d�w�5��������9��hY�*��h�4�
�:�$�����I�Ʃ�@�L�U���!�%�<�<�1��A܁�K���W�@��U¹�6��3�
�c��C������]��[��E���9�0�w�w�]�}�W���&����lR��h�I���d�u�=�;��0�(�������9��S�����;�!�9�f�`�}����[����V��U����