-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�c��m���}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e�'�3�4�'�<�G��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����T��U��������W�W���&ù��U9��G��E���
�9�u�u���3���>����F�G1�����4�%�4�d�m��W���&����p9��t:��U��u�:�;�:�g�f�W���	�֓�V ��[��*ۊ�%�#�1�o��}�#���6����9F���*���
�4�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���&����^��V�����u������4�ԜY�Ƽ�9��E��U���������!���6���F��@ ��U���_�u�u�
��8��������WF��~ ��!�����n�u�w�-�C�������T9��R1�Oʚ�������!���6���F��@ ��U���_�u�u�
�������֓�lV��G1����������4�ԜY�Ƽ�9��C�����
�
�u�u��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�M����Z��P1�����4�
�9�u�w��W���&����p]ǻN��*ފ�
�<�<�2�g�8�F��6����g"��x)��*�����}�d�3�*����P���F��1�����;�
�
�
��-����Cө��5��h"��<��u�u�%�a��)����&¹��F��x;��&���������W��Y����G	�UךU���
�
�
�<�>�:�F���H����E
��N��!ʆ�����]�}�W���&����Q��h^��U���������4���Y����W	��C��\�ߊu�u�
�
�2�����I����E
��N��U���
���n�w�}��������V��N�<����
�����#���Q����\��XN�N���u�%�`�'�1�?����&����_�'��&������_�w�}�(ف�&����]��h��U��� �u��
���(���-��� W��X����n�u�u�%�a���������V9��V�����u� �u����>��Y����lP��h�����d�0�e�o��	�$���5����l0��c!��]��1�"�!�u�~�W�W���&Ź��G��Y	��*���
�%�#�1�m��#ύ�=����z%��N������!�8�;���(���Y����`2��{!��6�����u�f�w�2����I��ƹF��hX��*���<�2�e�0�f�<�(���Y�ƃ�gF��s1��2���_�u�u�
�������ד�lW�!��U���
���
��	�%���Hӂ��]��G�U���%�c��!�:�3�(ށ�&¹��l��T�� ����
���l�}�WϮ�A����Z��P1����o������0���/����aF�N�����u�|�_�u�w��(�������lV��h^�����1�o�����;���:���F��1�����;�
�
�
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���YӖ��l%��^�����0�e�4�
�;�}�W���Y����)��tUךU���
�
�
�<�>�:�G���H����f2��c*��:���
�����l��������l�N��M���!�8�;�
���(������)��=��*����n�u�u�'�e�4�������9��N�:���������4���Y����W	��C��\�ߊu�u�
�
��4����H����l��A��Oʚ�������^�����Ɠ9��_�����0�7�=�#�8�}�Eٛ�O�ҍ�lV��DNךU���!�'�7�!�w��2���7����z)��~ ��U������_�w�}��������p)��h)��0�������w�;��������A��C�� ���<�_�u�u�:�k�4��8����[
��^��E���a�.��
���(���<΅��.��h'�� �����h�y���9���&����w[��"��<������h�4�'�E߽�����J��d1��%������g�y�m�G��1����}6��h/��=׺�=�'�y����(���:����S�� [�=�������d�q�;��� ����g[��Y��9����
��h�{��(���&����
J��d1��;���h�`�c����9���-�����=N��U���&�4�!�4��2��������F��d:��9����o�u�d�l�}�WϽ�����GF��h�����:�<�
�u�w�	�(���0����A��d��Uʶ�;�!�;�u�'��(���&����F��d:��9�������w�o��������\�^�W�ߊu�u�:�&�6�)����-����l ��h_��U���
���
��	�%���Y����G	�N�U��e�n�u�u�4�3����Y����g9��1����o������!���6�����Y��E���h�w�e�w�]�}�W���
������T�����f�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�u�W�W�������]��G1�����9�d�d�o���;���:����g)��^�����:�e�u�h�u��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�d�g�g�$���5����l0��c!��]���:�;�:�e�w�`�U���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�o�G��*����|!��h8��!���}�u�:�;�8�m�W��[���9F������!�4�
�:�$��݁�Y�Ɵ�w9��p'��#����u�d�1� �)�W���C���D��N�����!�;�u�%�4�3����K���5��h"��<������}�w�2����I����D��UװU���&�2�4�u�'��(���Y�Ɵ�w9��p'��#����u�g�1� �)�W���C���W�=N��U���'�7�!�u�$����������^ �����u�!�'�7�#�}��������]��QN��*���3�8�o�&�0�<�W���[����]ǻN�����9�4�
�<��.����&����U��N�&������_�w�}����Ӈ��@��U
��D���u����l�}�Wϭ�����C9��E�����4�e�<�
�>�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�����%�4�e�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���@��V��*ڊ�0�
�9�=����������@��N��1�����_�u�w�4����	�֓�V ��[��*ڊ�%�#�1�%�2�}�W���&����pF��I�N���u�&�2�4�w��(���&����R9��^ �����u��
����2���+������Y��E��u�u�&�2�6�}�(߁�����C��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�֓�V ��[��*ۊ�%�#�1�<��4�W���-����t/��=N��U���;�9�%�e�%�;�����ד�C9��S1�����u��
���}�J���^���F��P ��U���
�0�
�4��3����Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*ۊ�0�
�4�
�%�:�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��B�����Y�����'�3�8�-�6���������\��c*��:���n�u�u�&�0�<�W���&����^��V�����'�2�o����0���C���]ǻN�����9�%�g��%�2�(���
���5��h"��<������}�f�9� ���Y����F�D�����
�
�0�<�3�-����Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�D�����
�
�0�<�3�<�(���&����Z�=��*����n�u�u�$�:����&����A��h�����%�0�u�u���8���Y���A��N�����4�u�
�
�2�����I����@��N��1��������}�D�������V�=N��U���;�9�%�`�%�;����&ù��V�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�<�;�9�'�h��������9��h��*���&�2�o����0���s���@��V��*ߊ�0�
�0�4�g�<�(���&����\��c*��:���u�h�r�r�]�}�W�������lS��R�����d�<�
�<�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��E�����
�
�'�2�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�g�m�L���Yӕ��]��G1�����7�!�
�
�'�+����&����	F��s1��2���_�u�u�<�9�1��������V��1��*���
�'�2�o���;���:���V�=N��U���;�9�4�
�>�����K����q)��r/�����u�<�;�9�>���������C9��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:����5����u	��{��*Ҋ�
�0�
�`�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������C9��P1������&�g�3�:�l�Mύ�=����z%��N�����4�u�%�&�0�?���O����|)��v �U���&�2�4�u�:����I����	F��s1��2������u�g�9� ���Y����F�D�����8�
�0�
�a�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������C��ي� �f�m�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������`9��h(��*���%�g�
� �c�i����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*����'��:��n����L���5��h"��<������}�f�9� ���Y����F�D������9�
�:��2���&����W��N�&���������W��Y����G	�UךU���<�;�9�3��)�1���5����S��R	��M���u��
����2���+������Y��E��u�u�&�2�6�}�(ہ�&����]��B�����0�e�d�3��i�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����2�6�0�
��.�D������5��h"��<��u�u�&�2�6�}��������lW��T��:����n�u�u�$�:��������9��1��*��
�%�1�;�w�}�#���6����9F������%�a��!�:�3�(�������l��h\�� ��l�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����r9��Z��*���3�'�d�0�f�l����LŹ��\��c*��:���
�����l��������l�N�����u�
�
�
�>�4��������9��1�����c�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��l$��^�����3�0�
�
���(���M�֓� F��d:��9�������w�n�W������]ǻN�����9�%�c��#�0��������lW��h^��*���a�b�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��C����� �3�'�d�2�l�F���&����CU�=��*����
����u�FϺ�����O��N�����4�u�
�
��4��������A9��R1��G���
�l�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������l^��h�����7�3�0�
���(ށ�����l��N��1��������}�D�������V�=N��U���;�9�%�m��)����&����V��h��*؊� �`�`�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��t1�����
� �3�'�f�8�F�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�
����������U��1��D���3�
�d�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��*���
� �f�e�6�����Y�Ɵ�w9��p'�����u�<�;�9�0�-�����ד�F9��1��*���0�o�����4�ԜY�ƿ�T��	��*���
�
�
� �d�m��������	F��s1��2���_�u�u�<�9�1�����֓�lW��B1�E���
�0�
�9�?��W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����3�d�3�
�o���������lU�=��*����
����u�FϺ�����O��N�����4�u�'�
���(ށ�����l��g�����u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����U9��Q��Mڊ�;�'�3�7�#��W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����3�d�3�
�o���������F��d:��9�������w�n�W������]ǻN�����9�2�%�3�g�;�F���&����R��R����o������!���6���F��@ ��U���_�u�u�<�9�1�����֓�lW��B1�E���
�0� �;�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��*���
� �f�e�6��������5��h"��<������}�f�9� ���Y����F�D�����'�
�
�
�����I����A��E ��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���&����U��^�����!�'�
�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��1��D���
�m�
�%�4�}�W���&����p]ǻN�����9�%�c��#�0��������l��h_��*���
�d�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����q9��Z��*���3�'�0�d�g�.����K���5��h"��<������}�f�9� ���Y����F�D�����
�
�
�<�>�:��������9��D1����m�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�O����Z��P1�����
�
�
�
��8�(��Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y������!�8�;��(�����ד�l��R	��C���u��
����2���+������Y��E��u�u�&�2�6�}�(ہ�&����]��B�����d�e�&�'�0�o�@��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���<�<�2�7�1�8�(���&¹��A��W�Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�i�6�������Q��R��*ڊ�
�
�0�
�g�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�����;�
� �3�%�8�G���
����lU��T��!�����
����_������\F��d��Uʦ�2�4�u�
����������U��R1��D���'�2�f�l�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������l^��h�����7�3�0�
���(�������F��d:��9�������w�n�W������]ǻN�����9�%�m��#�0��������l��h_��*���
�`�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Z9��E1�����
�0�
�c�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������A��h^��*ۊ� �f�e�4��)����	����A��R	��U���
���u�j�z�P�ԜY�ƿ�T����;���&�u�u����>���<����N��S�����|�_�u�u�>�3�Ͽ�&����Q��\�Oʗ����_�w�}����Ӈ��@��U
��D��o�����W�W���������D�����f�u�u����L���Yӕ��]��V�����1�
�m�u�w��;���B�����Y�����<�
�1�
�a�g�5���<����F�D�����%�&�2�7�3�h�W���6����}]ǻN�����9�4�
�<��9�(��CӤ��#��d��Uʦ�2�4�u�%�$�:����A����q)��r/�����u�<�;�9�6���������\��x!��4��_�u�u�:�'�3����Kţ��R��h^��*����u�u�%�%�}�}���Y���R��[��U��������W�W���Y�ƭ�l��T��;ʆ�����]�}�W���Y����G��T��;ʆ�����]�}�W���Y����\��N��!ʆ�����]�}�W���Y����W
��N��!ʆ�����]�}�W���Y����V��T�� ����
���l�}�W���Yӏ��A��V����o��u����>���<����N��
�����e�n�u�u�w�}��������K9��N��U���
���
��	�%���Hӂ��]��G�U���u�u�<�
�2�4���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF�N�����3�7�!�
�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y���R��R����o������0���/����aF�N�����u�|�_�u�w�}�W�������]9��N��!ʆ�������8���J�ƨ�D��^����u�u�u�%�%�)����Y�ƃ�gF��s1��2������u�d�}�������9F�N��U���'�!�'�
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���Y�����E�����u�u� �u���8���&����|4�_�����:�e�n�u�w�}�WϿ�&����A��T�� ����
�����#���Q����\��XN�N���u�u�u�4��8�Mϗ�Y����)��tN����u�;�u�:�'�3���s���T��N�����3�e�3�d�1��O���Y����\��CN��C���m��
�
��W�W�������R�=N��U���u�%�6�>�j�}�������F�N��*���u�k�4�
�$�q�W���Y����C9��V��H���'�
�
�
�����I����@��CBךU���u�u�%�1�9�}�IϹ�	����l ��h��F���4�
�:�0�]�}�W���Y����W
��
P�����
�
�
�
�"�n�G���&����l�N��Uʴ�
�0�1�u�i�:����I����l ��V�����0�1�y�u�w�}�WϷ�&����R
��V1�H���'�
�
�
�����I����A��V����_�u�u�u�w�3��������[�P�����3�d�3�
�o���������lU�N��U���<�
�0�<�3�i�J�������9��1��*��
�;��'�8��[���Y�����E�����
�u�k�2�'�;�G���H���� ^��^ �����0�4�e�_�w�}�W���	����F��N��U���
�
�
�
��(�D�������G��h^�U���u�u�4�
�2�(���D�ƫ�C9��1��D���
�m�
�%�%�)����U���F������'�
�u�k�0�-�����ד�F9��1��*��� �;�g�_�w�}�W���	����F��N��U���
�
�
�
��(�D�������G��h]�U���u�u�4�
�2�(���D�ƫ�C9��1��D���
�m�
�%�%�)����U���F������'�
�u�k�0�-�����ד�F9��1��*��� �;�`�_�w�}�W���	����X��E��*ڊ�
�
� �f�g�<�(���B��Ɠ9l�N�U���u� �'�;�w�)��������l ��N��U���u�!�!�u�6�5���T���F��h-�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�6��$������R��c1��D���8�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�w�}�W���Y���F�N��U����
�&�u�j�<�(�������F�N��U���u�u�0�1�>�f�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�w�/�(���&����U��^�����4�!�4�
�#�/�(���Y����T��E�����x�_�u�u�%��(߁�&¹��lU��h�����!�4�
�!�%�����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��G1��E���d�3�
�m��-��������@��C1����u�%�6�;�#�1����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C\�����|�4�1�}�/�)����&����^��N�����:�&�
�#��t�^Ϫ���ƹF�N��U���u�u�u�u�%��(߁�&¹��lU��h�����!�4�
�!�%�����DӇ��P	��C1�����d�_�u�u�w�}�W���Y�Ʃ�@��F��*���&�
�:�<��}�W���&����U9��Q��Mڊ�%�'�4�,�~�)����Y���F�N��U���u�u�'�
���(ށ�����l��D�����
�!�'�
�2�}�JϿ�&����G9��P��E�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����lV��R�����
�
�%�#�3�-����
������T��[���_�u�u�
��8�(�������R��[
�����4�&�2�
�%�>�MϮ�������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�W��PӒ��]l�N��U���u�<�u�4��.�W���H����[��N��U���u�u�u�u�'�m��������lV��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�0�
�;�5�(߁�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������O��_�����u�u�u�u�w�}�W���Y���C9��E�����4�e�4�
�;�����E�Ƽ�9��Q1�����e�4�
�9�l�}�W���Y���F�N��U���u�3�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���
�9�=�
��/�Ͽ�
����C��R��U���u�u�%�e�%�;�����֓�A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�e�'�3�6�-����	����[��G1�����9�f�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʥ�e�'�3�4�'�<�G���&������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^�������9F�N��U���u�u�u�u�w��(���&����R9��G��U��%�e�'�3�6�-���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
��8�(�������R��[
�����4�&�2�u�%�>���T���F��1�����%�4�d�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���
�9�=�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���<�u�4�
�>�����A����[��=N��U���u�u�u�u�w�}�W���Y����A��V�����4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}�W���Y����_��F��*���
�1�
�c�w�5��ԜY���F�N��U���u�u�u�%�g�/����	����l��A�����u�h�%�e�%�;�����ד�C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(߁�����C��1�����&�<�;�%�8�8����T�����h��*���=�
�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l��h�����
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�m��������lW��G1�����u�=�;�_�w�}�W���Y���F�N��E���3�4�%�4�f�-����DӖ��l��h�����n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�����-�4�
�9��/�Ͽ�
����C��R��U���u�u�%�d�%�;��������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�2�����	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�<�(���&���� ^�����ߊu�u�u�u�w�}�W���Y���F��1�����-�4�
�9��/���Y����\��h�����n�u�u�u�w�}�W���Y�����^�����<�
�1�
�b�}����s���F�N��U���u�u�u�u�'�l��������C9��S1�����h�%�d�'�1�0����&����9F�N��U���u�u�u�u�w�3�W���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
��8�(���&������^	�����0�&�u�x�w�}��������R��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�d�%�;����	����[��G1�����9�f�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1�����-�4�
�9�~�t����Y���F�N��U���u�u�u�
��8�(���&����Z�G1�����8�-�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*���<�1�4�
�;���������]F��X�����x�u�u�%�e�����&����_��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�%�g��/����	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�<�(���&���� ^�����ߊu�u�u�u�w�}�W���Y���F��1�����
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W���Y���V
��QN�����2�7�1�c�~�)����Y���F�N��U���u�u�u�u����������E
��G��U��%�g��'�8��������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�g��%�2�(���Ӈ��Z��G�����u�x�u�u�'�o�'�������V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�0�<�3�-����DӇ��P	��C1��F؊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����c��X
�����1�|�u�=�9�W�W���Y���F�N��Uʥ�g��'�:��/���Y����c��X
�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����A��U��*ڊ�%�#�1�%�2�}����Ӗ��P��N����u�
�
�0��8��������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�2�����I����E
��G��U��4�
�:�&��2����B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�;�_���
����W��_�����u�u�u�u�w�}�W���Y���F���*���
�0�4�e�6��������F��h�����:�<�
�n�w�}�W���Y���F�N�����u�4�
�<��9�(��Y����l�N��U���u�u�u�u�w�}�WϮ�L����l��V1�����9�
�'�2�k�}�(ځ�����G��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����A��U��*ڊ�'�2�4�&�0�}����
���l�N��@���3�7�!�
��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h��*���4�e�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ځ�����G��h�����|�u�=�;�]�}�W���Y���F�N�����'�3�7�!������E�Ƽ�9��Q1�����n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�����!�
�
�%�!�9����Y����T��E�����x�_�u�u����������l��A�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(���&����lW��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�0�
�2�<�F���&����C��R�����:�&�
�:�>��L���Y���F�N��U���u�9�<�u�6���������F��R ��U���u�u�u�u�w�}�W���Y����lS��R�����d�4�
�9��/���Y����A��U��*ۊ�%�#�1�_�w�}�W���Y���F�N��ʼ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�����!�
�
�'�0�<����Y����V��C�U���%�`�'�3�5�)�(ށ�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ߊ�0�
�0�4�f�-����DӇ��P	��C1��F؊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����A��U��*ۊ�%�#�1�|�w�5��ԜY���F�N��U���u�%�`�'�1�?����&����Z�G1�����7�!�
�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����<��'��8��(���&����R��P �����&�{�x�_�w�}�;���&����	��hV�����c�
�&�<�9�-����Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�^�����<�
�1�
�`�t����Y���F�N��U���u�u�u��;���������l��h]�U��<�
�<��%�����&¹��T9��UךU���u�u�u�u�w�}����Yۇ��@��U
��D��u�=�;�_�w�}�W���Y���F�N��*����'��:������O�����T�����g�e�_�u�w�}�W���Y���V��^�U���u�u�u�u�2�9���s���F�R ����u�u�0�1�'�2����s���K�V�����'�6�&�{�z�W�W�������@F��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���^�Ƹ�VǻN��U���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o����H�ƭ�WF��O�����
� �f�m�'�}�W�������l
��h^��\ʡ�0�_�u�u�w�}�W���Y�ƪ�l
��q��9���
�f�'�2�b�m�K���*����u	��{��*���3�
�e�
�d�W�W���Y���F�N��*����'��:��h����L���F��h��3����:�
�`�1��Fށ�J���F�N��U���u�!�%�'�0�h�C��Y����U��^��D�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�E������F��R ךU���u�u�u�u�w�}�;���&����	��hV��*���
�`�u�h�>���������C9��1��*��
�g�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=N��U���4�&�2�u�%�>���T���F��X�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������A��N���ߊu�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�Փ�@��N��ʻ�!�}�%�6�9�)���������h��*���
� �f�e�6�����P����[��N��U���u�u�u�u�'�i�6�������Q��R��*ڊ�
�
�0�
�g�}�JϮ�M����Z��P1�����
�
�
�
��(�C���	��ƹF�N��U���u�u�
�
��4��������A9��1�����2�g�e�i�w��(�������l��Q��D���e�d�3�
�c��D�ԜY���F�N��Uʥ�a��!�8�9���������lV��h��*��u�h�%�a��)����&����V��h��*؊� �a�f�%�l�}�W���Y���F���*���<�<�2�7�1�8�(���&¹��A��X�I���
�
�
�<�>�:��������V9��1��*���
�f�_�u�w�}�W���Y���C9��u1�����
� �3�'�2�m�G�������W�
N��C���!�8�;�
�"�;�����֓�l ��Y����u�u�u�u�w�}�W���	�Г�l��^ �����0�
�
�
������J�����h,�����2�7�3�0���(߁�&����V��UךU���u�u�u�u�w�}�(ف�&����]��B�����d�e�&�'�0�o�B��Y����q9��Z��*���3�'�d�0�f�o����@¹��l�N��U���u�u�u�%�a���������U ��h��*ۊ�
�0�
�d�w�`����;����Z��U�����
�
�
�
�"�i�C���B���F�N��U���u�
�
�
�>�4��������V9��1�����f�c�i�u���(�������F ��E1�����d�3�
�l��n�}���Y���F�N������!�8�;��(�����֓�l��R	��G���h�%�m��#�0��������lW��h^��*���`�`�%�n�w�}�W���Y���F��hV��*���<�2�7�3�2��(ށ�&����T9��N�U���
�
�<�<�0�?����&¹��9��Q��D؊�f�_�u�u�w�}�W���Y�Ƽ�9��C����� �3�'�0�f�l��������Z�G1��6���8�;�
� �1�/�F���H�ԓ�F9��1��N���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B���F���U���!�&�4�0��-�9���
����UF��RN�����8�6�<�0�w�p�W�������l ��h�����%�:�u�u�%�>��������l ��N��*���u�%�&�2�5�9�F��Y����P	��1��*��
�g�u�'���(���&����V��G1�����u�u�7�2�9�}�W���YӅ��VF��h-�����<�_�u�u�w�}�W�������C9��h��*���
�u�k�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���&�2�7�1�f�i�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W���Y����_��N��U���u�u�u�u�w�}����*����Z�V��!���d�3�8�e�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����g9��1����h�u�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�1�
� �d�e����Y����\��h��*���|�u�=�;�w�}�W���Y���F�N�����
�&�u�h�6��#���H����lV��N��U���u�u�u�u�2�.�}���Y���F�N��U���4�
��3�:�a�W���*���� 9��Z1����u�u�u�u�w�}�W���Y����F�N��U���"�0�u�%���܁�
����X�N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������]��[����h�2�%�3�g�;�F���&����R��X ��\���!�0�_�u�w�}�W���Y���F�V��&���8�i�u�%���݁�
����9F�N��U���u�u�u�9�2�}�W���Y���F�N��U����
�&�u�j�<�(���
�Փ�@��d��U���u�u�u�u�w�8�Ϸ�B���F�N��U���;�:�=�'�w�c�W���Y���F�N��U����
�&�u�j��/���s���F�R �����n�u�u�0�3�-����
��ƹF�N��*���0�4�&�2�w�/����W���F�V�����4�&�2�
�%�>�MϮ�������T����<�
�&�$���݁�
������C��ي� �f�m�%�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�g�3�8�f�}��������K��X ��*���f�m�%�u�w�-��������lV�G�����_�u�u�u�w�}�W�������[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�:�2�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������]F��X�����x�u�u�4��9����
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�|�u�w�?����Y���F��QN�����}�%�6�;�#�1����H����C9��V��\ʴ�1�}�%�6�9�)���������D�����
��&�d�1�0�G���Y����l�N��U���u�4�
�1�2�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���'�4�,�4�$�:�W�������K��N�����0�1�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
�ԓ�@��N�����;�f�3�
�o��E�ԜY�Ʈ�T��N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!��.�(�������\�R�����f�3�
�m��o�JϿ�&����G9��1�\���!�0�u�u�w�}�W���YӇ��A��NN�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��h_�U���<�;�%�:�2�.�W��Y����C9��P1����a�4�&�2��/���	����@��G1�����u�
�
�0��1����&����_��Y1�����
�
�0�
�;�5�(ށ�	����l��D��U���
�0�
�4��-��������TJ��h\�����1�4�
�9��3����Y����A��U��*ڊ�%�#�1�<��4�[Ϯ�L����l��V1�����9�
�;�&�0�W�W�������F�N��U���u�u�4�
�>�����K���N��h\�����1�4�
�9��3����DӇ��P	��C1�����e�u�'�}����������l��h�����h�4�
�:�$�����&����AF��h[�����0�4�e�4��1�(���
�����T�����2�6�e�u�%�u�(ځ�����G��h�����<�
�<�u�w�-��������Z��N��U¥�e�'�3�4�'�<�G���&����Z��^	��U���6�;�!�9�0�>�G����μ�9��Q1�����d�4�
�9��3����DӇ��P	��C1�����e�u�'�}�'�.����DӇ��P	��C1�����e�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��o�W�������A	��D�X�ߊu�u�%�&�0�?���N����Z��G��U���'�6�&�}�'�.��������l��h��*���4�
�<�
�3��E���Y����V��=N��U���u�u�u�u�w�-��������Q�
N�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9��������T9��S1�A���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�a�w�.����	����@�CךU���%�&�2�7�3�l�A���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z������!�9�d�d�j�<�(��������Y��D���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�c�w�.����	����@�CךU���%�&�2�7�3�l�A���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������Z������!�9�d�d�j�<�(��������Y��G���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�b�w�.����	����@�CךU���%�&�2�7�3�l�E���
����C��T�����&�}�%�&�0�>����-����l ��h\����3�e�3�d�1��O߁�	����VOǻN�����_�u�u�u�w�}�W���Y����Z��S
��B���h�}�4�
�8�.�(�������F��h��*���$��
�!��.�(�������\�V�����
�:�<�
�w�}����&ù��9��h]�*���1�;�|�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(������]F��X�����x�u�u�4��4�(���&�ߓ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��N�U´�
��3�8�g�9� ���Y�����T�����d�d�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�n�W�������A	��D�X�ߊu�u�%�&�0�?���&����T��E��Oʥ�:�0�&�4��)�������T9��R��!���d�3�8�e�w��(���&����R9��V�����u�u�7�2�9�}�W���Y���F������7�1�f�u�j�u��������_	��T1�Hʥ�e�'�3�4�'�<�G���&������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^��Y����]��E����_�u�u�x�w�-��������W��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��V�����2�
�'�6�m�-����
ۇ��@��T��*���&�g�3�8�f�}��������U��V��G�ߊu�u�0�<�]�}�W���Y���F�V�����1�
�m�u�j�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����0�<�6�;�d�;�(��&�����T�����d�e�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�C���
������T��[���_�u�u�%�$�:����MŹ��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(߁�����C��1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�a�w�`�_���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����u�;�u�4��2��������F�G1�����4�%�4�d�6�����B����������n�_�u�u�z�}��������lS��V�����'�6�&�{�z�W�W���	����l��h[�����2�
�'�6�m�-����
ۇ��@��CB�����2�6�0�
��.�F������C9��E�����4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�B���D�΢�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�d�'�3�8�/�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��N�����u�'�6�&�y�p�}���Y����Z��S
��A���&�2�
�'�4�g��������C9��V��U���&�2�6�0��	��������F��1�����
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�0�<�3�<�(���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��N�����u�'�6�&�y�p�}���Y����Z��S
��D���&�2�
�'�4�g��������C9��V��U���&�2�6�0��	��������F��1�����!�
�
�%�!�9�}���Y����]l�N��U���u�u�u�4��4�(���&���F��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
�2�����I����E
��UךU���;�u�'�6�$�f�}���Y���R��^	�����e�4�&�2�w�/����W���F�V�����1�
�e�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�`�'�3�7�#��(������F�U�����u�u�u�u�w�}�WϿ�&����Q��^��H���:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ځ�����G��h�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���ށ�
����R��P �����&�{�x�_�w�}��������B9��h��*���
�
�&�<�9�-����Y����V��V�����1�
�l�_�w�}����s���F�^�����<�
�1�
�n�}����s���F�N�����<�
�&�$���ށ�
����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����U��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�V�����&�$��
�#�����Y����T��E�����x�_�u�u�'�.��������l��h��*ۊ�&�<�;�%�8�}�W�������R��^	�����a�|�u�u�5�:����Y����������7�1�d�c�w�5��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�d�_�w�}�W������F�N��U���4�
�<�
�$�,�$�������^9��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h��*���$��
�!��.�(���
������T��[���_�u�u�%�$�:����&����GU��D��*���<�;�%�:�w�}����
�έ�l��h��*��|�u�u�7�0�3�W���Y����UF��G1�����1�d�c�u�?�3�}���Y���F�V�����&�$��
�#�����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�<�
�&�&��(���&����F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����P	��1��*��
�g�i�u�f�}����Q����Z9��E1�����
�0�
�c�w�}��������ET��N�����e�n�u�u�1���������C9��h��A���%�u�h�_�w�}�W���&ù��U9��G��D���
�<�u�=�9�u��������l��G��U��|�0�&�u�w�}�W���	�֓�V ��[��*ڊ�;�&�2�_�w�}�$���&����	��h\�����d�
�f�i�w�}�W���YӖ��l��h�����<�
�<�u�?�3�_���&����V��F�U���d�|�0�&�w�}�W���YӖ��l��h�����<�
�<�n�]�}�W������lV��h_�� ��e�4�
�0�6�.��������@H�d��Uʲ�%�3�e�3�f�;�(��&����V9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�
�&��q��������l ��V�����4�
�<�
�$�,�$�������^9��=N��U���<�_�u�u�w�}����Q����\��h�����u�u�%�6�~�<��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����P	��1��*��
�g�h�4��2����¹��O����ߊu�u�u�u�w�}����&ù��9��h]�*���6�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����U9��Q1�����m�
�%�6�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߊu�u�'�
���(ށ�����l��D����u�'�
�
���(���J�֓�C9��V�����!�'�
�0�l�}�WϹ�	����l ��h��F���<�
�0�<�3�i�K���&����A��h�����_�u�u�'���(���&����V��Y1�����%�4�d�i�w���������\��1�����e�_�u�u�%��(߁�&¹��lU��h�����7�!�
�u�j�;�(���?����\	��[�����m�n�u�u�0�-�����ד�F9��1��*���
�4�
�u�j�-�F�������l��D�����u��9�
�8�����A�ד�F9��1��U��&�1�9�2�4�+����Q����T�������:�
�:�%�o�/���A���F��P ��]���6�;�!�9�e�l�^�ԶY���F��1�����%�4�e�4��1�(���
����@��YN�����&�u�x�u�w�-�G�������[��h�����<�
�<�
�$�4��������C��R�����'�3�4�%�6�m��������lV��R�����
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1�����4�%�4�e�6�����Y����l�N��U���u�%�e�'�1�<����I����E
��^ �����h�%�e�'�1�<����I����E
��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��Q1�����e�4�
�9��3����E�Ƽ�9��Q1�����e�4�
�9��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�G1�����4�%�4�e�>�����
������T��[���_�u�u�
��8�(�������Z��^	�����;�%�:�u�w�/����Q����A��V����u�
�
�0��1����&����F��1�����%�4�e�4��1�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��1�����%�4�e�4��1�^������F�N��U���%�e�'�3�6�-��������TF���*���
�9�=�
�l�}�W���YӃ��VFǻN��U���u�u�
�
�2�����&ù��l��R�����'�3�4�%�6�m����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ڊ�0�
�9�=����������@��V�����'�6�&�{�z�W�W���&ù��U9��G��D���
�9�
�;�$�:��������\������}�
�
�0��1����&����_�G1�����4�%�4�d�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�0�
�9�?��(��������YNךU���u�u�u�u����������9��h��*���&�2�i�u����������9��h��N���u�u�u�0�$�}�W���Y���F��h^�����9�=�
�
�'�+����&����[��h^�����9�=�
�
�'�+������ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�0�
�9�?��(���
����@��YN�����&�u�x�u�w�-�G�������[��h�����4�&�2�
�%�>�MϮ�������h��*���=�
�y�%�g�/����	����l��PB��*ڊ�0�
�9�=���������F��P��U���u�u�<�u��-��������Z��S��*ڊ�0�
�9�=����������[��=N��U���u�u�u�
��8�(�������Z��^	��Hʥ�e�'�3�4�'�<�F�ԜY���F��D��U���u�u�u�u�'�m��������lW��Y1����u�
�
�0��1����&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�d�'�3�:�%��������l�������%�:�0�&�w�p�W���	�ד�V ��V�����1�<�
�<��.����	����	F��X��¥�d�'�3�8�/�<�(���UӖ��l��h��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��Q1�����
�9�|�u�?�3�}���Y���F�G1�����8�-�4�
�;��������C9��E�����4�
�9�n�w�}�W�������9F�N��U���u�
�
�0��<�(�������]9��PN�U���
�0�
�4��-����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�0�
�6�����Ӈ��Z��G�����u�x�u�u�'�l��������]9��P1�����
�'�6�o�'�2����	�ד�V ��V����'�3�8�-�'�8�[Ϯ�H����l��h�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�F�������l��A��\ʡ�0�u�u�u�w�}�W���	�ד�V ��V�����2�i�u�
��8�(���B���F����ߊu�u�u�u�w�}�(ށ�����K9��h��U��%�d�'�3�:�%����B���F���U���u�u�u�0�3�-����
��ƓF�C��*؊�0�<�1�4��1�(���
����@��YN�����&�u�x�u�w�-�E�������R��[
�����2�4�&�2��/���	����@��h\�����1�4�
�9�{�-�E�������R��[
�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�E�������R��[
��U���;�_�u�u�w�}�W���&����A��h�����<�
�<�u�j�-�E�������R��[
�U���u�u�0�&�w�}�W���Y�����h>�����4�
�9�
�9�.���Y����c��X
�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l6��^�����<�u�&�<�9�-����
���9F���*���<�1�<�
�>���������PF��G�����%�g��'�8�q����)����W9��R	�����'�:�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h\�����1�4�
�9�~�}����s���F�N������'�:�
�9�.���Y����c��X
�U���u�u�0�&�w�}�W���Y�����h>�����<�
�<�u�j�-�E�������C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���%�a��!�:�3�(߁�&�����h/�����2�7�3�0���(߁�&���� V��=d��U���u�
�
�
�>�4�����֓�C9��SN�����u�'�6�&�y�p�}���Y����r9��Z��*ڊ�
�
�%�#�3�<����&����\��E�����%�6�y�4��4�(�������@��Q��D���-�!�:�1��(�D���	��ƹF��R	�����u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�E������R��Y��]���!�:�1�
�"�n�O���Y�ƭ�l��D��ۊ�|�|�u�=�9�W�W���Y���F��1�����;�
�
�
��-����E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���
�
�<�<�0�m��������WF������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����r9��Z��*ڊ�
�u�h�%�c���������U ��h��*ڊ�
�0�
�b�l�W�W���TӖ��l'��^�����0�d�4�
�;�}����Ӗ��P��N����u�
�
�
�>�4�����ד�C9��S1�����
�'�6�o�'�2��������F��h��*���$��
�!��.�(������\��h��F���%�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��G���8�d�u�;�w�2�_ǻ�����WU��B1�M���u�u�%�6�9�)����I�����YNךU���u�u�u�u���(�������l��h�����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϮ�M����Z��P1�����4�
�9�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�
�
�
�>�4�������F��1�����;�
� �3�%�8�G���
����lT��dךU���x�%�a��#�0����&����R��[
�����;�%�:�0�$�}�Z���YӖ��l'��^�����0�e�4�
�;���������PF��G�����4�
�0�u�'�.��������l��h��*���0�<�6�;�d�;�(��&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���݁�
������ ��]°�<�6�;�f�1��Oׁ�K����C9��Y�����e�|�|�!�2�}�W���Y���F��hZ��*���<�2�d�0�g�<�(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʥ�a��!�8�9��(���&����_�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}���YӖ��l'��^�����0�d�i�u���(�������F ��E1��D���&�'�2�g�c�W�W���T�Ƽ�9��C�����
�
�
�%�!�9�����Ƽ�\��D@��X���u�%�a��#�0����&����R��[
�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�e�;���Y����P	��1��*��
�g�_�u�w�8��ԜY���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��؊�&�
�|�4�3�3��������]��Q��MҊ�g�h�4�
�8�.�(���&���F��R ��U���u�u�u�u�'�i�6�������9��1��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���&ǹ��G��Y	��*���
�%�#�1�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R�����u�%�a��#�0��������lW��h^��*���a�g�%�u�j�W�W���Y�ƫ�C9��1��D���
�m�
�%�%�)����Y����N��G1�����a�e�u�u�f�t����Y���F���*���<�<�2�7�1�8�(���&¹��A��W����u�
�
�
�>�4��������9��1�����a�
�f�i�w�}�W���YӖ��l'��^�����3�0�
�
���(���&����D��F�����2�`�a�e�w�}�F�������9F�N��U���
�
�
�
��(�D�������G��h^�U���%�a��!�:�3�(�������l��h_�� ��c�%�u�h�]�}�W���Y����U9��Q1�����m�
�%�'�#�/�(������G��E��@��e�u�u�d�~�8����Y���F��hZ��*���<�2�7�3�2��(ށ�&����T9��UךU���
�
�
�<�>�:��������V9��1��*��
�f�i�u�w�}�W���	�ғ�l��^ �����0�
�
�
������N�ƻ�V�C�����`�a�e�u�w�l�^ϻ�
��ƹF�N�����
�
�
�
�"�n�G���&����A��dךU���x�%�`�'�1�?����&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��E�����
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�b�/��������R��[
����'�3�7�!����������TOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�`�'�3�5�)�(߁�	����O��_�����u�u�u�u�w��(���&����lV��G1�����
�<�u�h�'�h��������9��h��N���u�u�u�0�$�}�W���Y���F��h[�����0�4�e�4��1�(���
���F��1�����!�
�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ߊ�0�
�0�4�g�4�(���Y����T��E�����x�_�u�u����������l��D�����2�
�'�6�m�-����
ۖ��l��h����u�
�
�0��8����	������h��*���4�e�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��E�����
�
�%�#�3�t����Y���F�N��U���
�0�
�0�6�m���������h��*���4�e�_�u�w�}�W������F�N��Uʥ�`�'�3�7�#��(���
���F��1�����!�
�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��E�����
�
�%�#�3�4�(���Y����T��E�����x�_�u�u����������l��A�����<�
�&�<�9�-����Y����V��G1�����7�!�
�
�'�+����&ƹ��U9��C��*���#�1�%�0�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��Q1�����
�%�#�1�~�)����Y���F�N��*ߊ�0�
�0�4�f�<�(���&����Z�
N��@���3�7�!�
��-����s���F�R��U���u�u�u�u�w�-�B�������R9��V�����;�&�2�i�w��(���&����lW��G1�����0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�L����l��V1�����<�u�&�<�9�-����
���9F���*���
�0�4�d�>�����
����l��TN����0�&�%�`�%�;����&����lS��R�����d�%�0�y�'�h��������9��h��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u����������l��A��\ʡ�0�u�u�u�w�}�W���	�ӓ�V ��R��D���
�<�u�h�'�h��������]ǻN��U���9�0�_�u�w�}�W���Y����A��U��*ۊ�;�&�2�i�w��(���&����lW��E�����u�u�u�;�w�;�W���YӃ����T��N�ߊu�u�
�
��4����I����Z�G1��7���8�;�
� �1�/����I����V��_����u�x�%�c��)����&ù��9��h��U���<�;�%�:�2�.�W��Y����lP��h�����e�0�e�4��1�(�������A	��N�����&�4�
�0�w�-��������`2��C\�����y�0�<�6�9�n����A˹��l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����0�<�6�;�d�;�(��&�����T�����d�e�|�|�#�8�W���Y���F���*���<�<�2�e�2�m���������T�����2�6�d�_�w�}�W������F�N��U���%�c��!�:�3�(߁�&ù��l��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��ԶY����lP��h�����e�0�d�i�w��(�������l��Q�����e�&�'�2�e�h�}���Y���C9��u1�����
�
�
�
�'�+�Ͽ�
����C��R��U���u�u�%�c��)����&ù��9��h��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�o����H�Ʃ�Z��Y
�����m�
�g�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9����Q����P	��1��*��
�g�h�4��2����¹��O�C��U���u�u�u�u�w�-�A�������T9��R1�����9�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����q9��Z��*ڊ�
�
�%�#�3�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠu�u�%�c��)����&¹��F���*���<�<�2�7�1�8�(���&¹��A��]����u�x�u�
�������ד�lV��G1��ʴ�&�2�u�'�4�.�Y��s���C9��u1�����
�
�
�
�'�+����
����C��T�����&�}�%�6�{�<�(���&����l5��D�����d�u�-�!�8�9�(���J�ޓ�OǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���K����lW�V �����}�-�!�:�3����A����F��h�����#�
�|�|�w�5��ԜY���F�N��C���!�8�;�
���(������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�
�
�
�>�4�����֓�C9��SN�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���C9��u1�����
�
�
�u�j�-�A�������T9��Q��*���
�
�
�0��l�L�ԜY�����h,�����2�d�0�d�6�����
������T��[���_�u�u�
�������ד�lW��G1�����&�2�
�'�4�g��������C9��N��*���
�&�$���)�(���&����K��X ��*���f�m�%�|�w�}�������F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���g�3�8�d�w�3�W���Qۃ��G��S]�� ��m�%�u�u�'�>�����ד�O����ߊu�u�u�u�w�}�(ف�&����]��h��*���#�1�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӖ��l$��^�����0�d�4�
�;�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�
����������U��1��E���3�
�b�
�d�a�W���Y�����h��*���
� �f�e�6���������[����*���
�c�}�|�j�z�P������F�N������!�8�;��(�����֓�l��R	��F��u�u�%�c��)����&����V��h��*؊� �a�b�%�w�`�}���Y���C9��u1�����
� �3�'�2�m�G�������W��_��]���
�0�
�c��t�J���^�Ʃ�@�N��U���2�%�3�e�1�l����Aù��l��B��G�ߊu�u�
�
��4��������A9��R1��D���
�m�
�f�k�}�W���Y����A��h^��*ۊ� �f�e�4��8����Jӑ��]F��Z�����c�}�|�h�p�z�W������F�N��C���!�8�;�
�"�;����H�ד�l��h\�N���u�%�c��#�0��������lW��h_��*���a�d�%�u�j�W�W���Y�Ƽ�9��C����� �3�'�0�f�m����������YN�����0�
�c�}�~�`�P���Y����l�N��Uʲ�%�3�e�3�f�;�(��&����V��Y1����u�
�
�
�>�4�������F��1�����;�
� �3�%�8�G���
����lU��dךU���x�%�m��#�0����&����R��[
�����;�%�:�0�$�}�Z���YӖ��l%��^�����0�e�4�
�;���������PF��G�����4�
�0�u�'�.��������l��h��*���0�<�6�;�d�;�(��&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���݁�
������ ��]°�<�6�;�f�1��Oׁ�K����C9��Y�����e�|�|�!�2�}�W���Y���F��hV��*���<�2�e�0�g�<�(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʥ�m��!�8�9��(���&����_�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}���YӖ��l%��^�����0�d�i�u���(�������F ��E1��D���&�'�2�f�e�W�W���T�Ƽ�9��C�����
�
�
�%�!�9�����Ƽ�\��D@��X���u�%�m��#�0����&����R��[
�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�e�;���Y����P	��1��*��
�g�_�u�w�8��ԜY���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��؊�&�
�|�4�3�3��������]��Q��MҊ�g�h�4�
�8�.�(���&���F��R ��U���u�u�u�u�'�e�4�������9��1��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���&˹��G��Y	��*���
�%�#�1�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R�����u�%�m��#�0����&����[��hV��*���<�2�7�3�2��(߁�&����T9��UװU���x�u�
�
��4����H����l��A�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��C�����
�
�
�%�!�9��������\������}�%�6�y�6�����
����g9��1����u�-�!�:�3����A����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������F��SN�����-�!�:�1��(�D���	���R��X ��*���
�|�|�u�?�3�}���Y���F�G1��6���8�;�
�
���������R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���
�
�
�<�>�:�F���I����E
��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԜY�Ƽ�9��C�����
�
�u�h�'�e�4�������Q��R��*ۊ�
�
�0�
�b�f�}���Y����l^��h�����d�0�d�4��1�W�������A	��D�X�ߊu�u�
�
��4����H����l��A�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�����UӃ��G��S]�� ��m�%�|�u�w�?����Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�d�u�9�}��������\��h��F���%�u�u�%�4�3����H���O��_�����u�u�u�u�w��(�������lW��h_�����1�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W���	�ޓ�l��^ ��D���d�4�
�9�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߊu�u�
�
��4��������A9��R1��D���
�l�
�f�k�}�W���Y����l^��h�����7�3�0�
���(�������F��R �����'�2�`�a�g�}�W��PӃ��VFǻN��U���'�
�
�
�����I����A��E ��N���u�%�m��#�0��������lW��h^��*���`�`�%�u�j�W�W���Y�ƫ�C9��1��D���
�m�
�%�%�)����Y����N��G1�����a�e�u�u�f�t����Y���F���*���<�<�2�7�1�8�(���&¹��A��\����u�
�
�
�>�4��������9��1�����d�
�f�i�w�}�W���YӖ��l%��^�����3�0�
�
���(���&����D��F�����2�`�a�e�w�}�F�������9F�N��U���
�
�
�
��(�D�������G��h[�U���%�m��!�:�3�(�������l��h\�� ���l�%�u�h�]�}�W���Y����U9��Q1�����m�
�%�'�#�/�(������G��E��@��e�u�u�d�~�8����Y���F��hV��*���<�2�7�3�2��(ށ�&����T9��UךU���8�
� �a�g�-�W������l ��h"�����'�2�f�m�f�p�FϺ�����O��R �����#�_