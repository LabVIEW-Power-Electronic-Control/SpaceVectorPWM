-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�m�m�d�a���(���
����GF�N�����9�u�u����;���:���F��h��U���������}���Y����G��T��;ʆ�����]�}�W�������	F��cN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�%�<���6����g"��x)��N���u�<�
�%�%�8���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF��Y1�����
�u�u����;���:����g)��]����!�u�|�_�w�}��������G9��N��U���
���
��	�%���Hӂ��]��G�U���<�
�%�'�2�)�E��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����E�����u�u� �u���8���&����|4�_�����:�e�n�u�w�<�(�������\��b:��!�����
����_������\F��d��Uʴ�
�0� �;�e�g�8���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƭ�l��B��F��������4���:����U��S�����|�_�u�u�'�/����&����|3��d:��9�������w�n�W������]ǻN�����!�'�
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W�������\��yN��1�����|�_�9�f�}������P��RN�����:�u���f���������@FǻN�����4�!�4�
�8�.�(�������	F��s1��2���o�u�d�n�w�}��������R��X ��*���<�
�u�u���8���Y���A��N�����!�;�u�%���ށ�
����	F��s1��2������u�b�9� ���Y���F�^�D��u�u�6�;�#�3�W���*����9��Z1�Oʆ�������8���Lӂ��]��G��H���e�e�e�n�w�}��������R��c1��F���8�g�o����0���/����aF�
�����e�u�h�w�g�l�G��Y����\��V ������&�a�3�:�n�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���I����]ǻN�����4�!�4�
��.�B������5��h"��<������}�w�2����I����D��^�W�ߊu�u�:�&�6�)����-����l ��h[��U���
���
��	�%���Y����G	�N�U��e�e�w�_�w�}��������C9��Y����
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�e�w�]�}�W���
������T�����d�d�o����0���/����aF�
�����e�u�h�w�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�l�U�ԜY�Ư�]��Y�����;�!�9�d�g�g�$���5����l0��c!��]���:�;�:�e�w�`�U���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)����I����g"��x)��*�����}�u�8�3���Y���V�=N��U���&�4�!�4��2��������	F��s1��2������u�f�9� ���Y���F�L�U���6�;�!�;�w�-��������lW�=��*����
����u�W������F��L�W�ߊu�u�:�&�6�)��������_��h]��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��_�D��n�u�u�6�9�)����	����@��A]��F���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�D��e�w�_�u�w�2����Ӈ��P	��C1��F؊��o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��d�d�e�n�w�}��������R��X ��*���f�e�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�n�w�}��������R��X ��*���g�a�f�o���;���:����g)��_����!�u�|�o�w�m�G��H����D��N�����!�;�u�%�4�3����H¹�� F��d:��9�������w�l�W������F��L�E��d�e�d�n�w�}��������R��X ��*���g��o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�d�l�}�WϽ�����GF��h�����#�d�e�o���;���:����g)��_����!�u�|�o�w�m�G��I����]ǻN�����4�!�4�
�8�.�(���K����\��c*��:���
�����l��������\�_�D��d�d�e�n�w�}��������R��X ��*���g�f�u�u���8���&����|4�_�����:�e�u�h�u�m�G��H����]ǻN�����4�!�4�
�8�.�(���&����`2��{!��6�����u�`�3�*����P���V��^�N���u�6�;�!�9�}��������EP��N�&���������W������\F��T��W��d�e�n�u�w�>�����ƭ�l��D�����e�o�����4���:����S��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
����T��T��!�����
����_������\F��T��W��e�e�e�e�g�f�W�������R��V�����
�#�g�f�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����W��UךU���:�&�4�!�6�����&����F��d:��9�������w�k��������\�^�E��w�_�u�u�8�.��������]��[�*������o���;���:����g)��]����!�u�|�o�w�l�F��H����W��_�D��d�d�d�d�f�f�W�������R��V�����
�#�g���g�$���5����l0��c!��]��1�"�!�u�~�g�W��H����W��L�U���6�;�!�;�w�-��������9��q(��3�����u�u���8���&����|4�]�����:�e�u�h�u�l�F��H����W��_�D��d�d�d�d�f�l�F��H����W��_�D��u�u�6�;�#�3�W�������l
��1��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�D��w�_�u�u�8�.��������]��[�*��o������!���6���F��@ ��U���o�u�e�e�g�l�G��[���F��Y�����%�6�;�!�;�l�(��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��_�E��n�_�u�u�>�3�Ͽ�&����@�=��*����
����u�W������F��L�E��w�_�u�u�#�/����Y����V��S��U���!�<�2�_�w�}��������U��R �����u�3�4�
��;���
����_F��L�����_�u�u�<�9�1��������V��c1��D���8�e�o����0���s���@��V�����2�7�1�g�w�}�8���8��ƹF��^	��ʴ�
�<�
�&�&��(���&����F��d:��9����_�u�u�>�3�Ͽ�&����Q��V��U�����n�u�w�.����Y����U��\��D��������4���Y����W	��C��\�ߊu�u�<�;�;�;�(�������^9��h��*��a�o�����4���:����U��S�����|�_�u�u�>�3�Ϸ�&����\��X��Dۊ� �g�e�%�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������9��h(��*���%�d�
�0��l�E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V�����&�$��
�#�����Y�Ɵ�w9��p'�����u�<�;�9�6���������\��x!��4��u�u�&�2�6�}��������lT��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2���������Q�=��*����
����u�W������]ǻN�����9�0�<�6�9����M����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�g�1��Bׁ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�
�0��l�B��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��Q=��8���,� �
�f�1��Fׁ�K����g"��x)��*�����}�d�3�*����P���F��P ��U���-� ���#�o�(���&����\��c*��:���
�����l��������l�N�����u�&�0�
�2��F��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*���
�&�$���)�(���&����`2��{!��6�ߊu�u�<�;�;�<�(���&����
R�,��9���n�u�u�&�0�<�W���&�Փ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������_��N��1��������}�B�������V�=N��U���;�9�!�%�f����K����	F��s1��2������u�g�9� ���Y����F�D�����8�
�l�'�0�l�N���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��(�����a�
�g�o���;���:����g)��_����!�u�|�_�w�}����Ӡ��A��\�U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_�������V�=N��U���;�9�!�%�e�����K���5��h"��<������}�w�2����I��ƹF��^	��ʼ�8�b�3�
�`��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��^��B���2�d�d�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lP��Q��LҊ�f�o�����4���:����S��X����n�u�u�&�0�<�W���&�֓�V��\�Oʆ�������8���Lӂ��]��G�U���&�2�4�u��<�E�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�
�6�o�B�������
F��d:��9�������w�n�W������]ǻN�����9�4�
�<��.����&����U��N�&������_�w�}����Ӈ��@��U
��D��o�����W�W���������D�����'�2�d�f�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������l��h_�E��������4���Y����\��XN�N���u�&�2�4�w�8����&����@9��hW�*��o������!���6�����Y��E��u�u�&�2�6�}��������A	��E��D��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1�%���¹��_9��R��*���m�3�
�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��Y	��*���
�;�&�g�>�l�(���&����\��c*��:���
�����}�������9F������4�'�9�
�8�����Hʹ��V9��1��*��c�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Z��D��&���!�
�&�
�w�}�#���6����9F������4�
�<�
�3��D���Y����v'��=N��U���;�9�4�'�;���������
9��R1��F���
�e�e�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����R��[�����:�%�d�
���(ځ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�'��)�1���5����_��h��*ۊ� �d�m�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��3����:�
�l�e�8�F�������
^��N�&���������W��Y����G	�UךU���<�;�9�4�%�1�(���&����lW��1��D���3�
�d�g�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h'��0����0�8�a���(���&����	F��s1��2������u�d�}�������9F������6�
��������Mǹ��9��P1�C��������4���Y����W	��C��\�ߊu�u�<�;�;�<����&����	��h_��G���e�c�'�2�f�e�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�����'��:�
�n�o��������V�=��*����
����u�FϺ�����O��N�����4�u�9����%�������l��h��*��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���0����r4��R��A܊�
�
�0�
�n�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��3����:�
�
�2��G���Y����)��t1��6���u�d�1�"�#�}�^�ԜY�ƿ�T���������!�g��(�E���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�
���,�"��D���&����CW�=��*����
����u�FϺ�����O��N�����4�u�'�
�"�o�E���Y�Ɵ�w9��p'��#����u�c�u�8�3���B�����Y�����&�2�
� �e�h����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����%�
� �g�e�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��S1�����
� �g�`�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��R	��*���f�m�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ʃ�C9��G1�����g�
�a�o���;���:����g)��_����!�u�|�_�w�}����Ӓ��lR��Q��D؊�d�o�����4���:����P��S�����|�_�u�u�>�3�Ϫ�	����F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��n����NŹ��\��c*��:���
�����l��������l�N�����u�8�
�l�1��Oׁ�H����g"��x)��*�����}�u�8�3���B�����Y�����f�
� �f�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h�����l�
�g�o���;���:����g)��[�����:�e�n�u�w�.����Y����^��B1�C���u�u��
���(���-���T��X����n�u�u�&�0�<�W�������lW��Q��Dي�d�o�����4���:����S��S�����|�_�u�u�>�3�ϳ�����l ��_�����u��
����2���+������Y��E��u�u�&�2�6�}����I����U��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�o�(���M�ӓ�F��d:��9�������w�l�W������]ǻN�����9��
�
�"�i�G���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y������3�
�g��n�Mύ�=����z%��r-��'���f�1�"�!�w�t�}���Y����R
��Z��@���
�c�
�a�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��h��A���%�u�u����>���<����N��
�����e�n�u�u�$�:����K�ԓ�R��Q��A݊�d�o�����4���:����U��S�����|�_�u�u�>�3�Ϸ�����lR��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��A���&����CT�=��*����
����u�FϺ�����O��N�����4�u�8�
�`�;�(��&���5��h"��<������}�d�9� ���Y����F�D�����8�
�m�3��d�(��Cӵ��l*��~-��0����}�f�1� �)�W���s���@��V�����a�3�
�`��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���`�d�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƿ�\��R��*���`�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��@���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l��C1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������9��h[�*��o������!���6�����Y��E��u�u�&�2�6�}����N����U��G]��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�k�(���L�ߓ�F��d:��9�������w�h�W������]ǻN�����9�!�%�c��(�B���	����`2��{!��6�����u�`�w�2����I��ƹF��^	��ʡ�%�c�
� �b�e����Y����)��t1��6���u�`�u�:�9�2�G��Y����Z��[N��'���9�
�
� �b�i����Y����)��t1��6���u�`�u�:�9�2�G��Y����Z��[N����
� �`�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������V��F���
�d�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������^��1��*��
�d�o����0���/����aF�
�����e�n�u�u�$�:����&����P��N�&���������W������\F��d��Uʦ�2�4�u�
�����J����	F��s1��2������u�g�9� ���Y����F�D�����7�3�
�a��n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h�����d�3�
�l��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���c�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�e��hZ�� ��l�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Q��B1�@���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Oƹ��lS��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2���������9��T��!�����
����_�������V�=N��U���;�9�!�%�1��Cށ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�e�3��i�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�
� �c�n�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��D�����a�1�8�'�6����H����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�d��(�A���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʦ�:�0�0�2�����J����	F��s1��2������u�d�}�������9F������!�%�f�
�"�k�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����3�
�m�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������
9��hY�*��o������!���6�����Y��E��u�u�&�2�6�}��������U��[��D��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����P��N�&���������W��Y����G	�UךU���<�;�9�!�'�i�(���N�֓�F��d:��9�������w�h�W������]ǻN�����9�9�
� �`�k����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���b�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ�� T��B1�E���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����N¹��lQ��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��C���&����CT�=��*����
����u�W������]ǻN�����9�'�#�
�"�j�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����6�&�
� �a�i����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N����
� �b�m�'�}�W���&����p9��t:��U���u�:�;�:�g�f�W���
����_F��Y	��*���
� �b�g�'�}�W���&����p9��t:��U���u�:�;�:�g�f�W���
����_F��a1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������]��h�� ��g�%�u�u���8���&����|4�N�����u�|�_�u�w�4����+����9��[1����� �b�a�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������R��1�����0�
�
�
�"�e�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����d�4�9�:�2��(���N�Г�F��d:��9�������w�m��������l�N�����u�8�
�c�1��E߁�K����g"��x)��*�����}�u�8�3���B�����Y��'���0�
�9�
�2�2�(���A�Г�F��d:��9�������w�m��������l�N�����u�4�2�d�6�1����
�ד�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Cہ�����l^��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��O���&����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�n����O����\��c*��:���
�����}�������9F������&�9�!�%�c�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʺ�
�:�1�f�>�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʇ�;�0�
�9��3����&����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�h����Nǹ��\��c*��:���
�����}�������9F������%�l�
�
�"�e�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V��*���<�3�
�f��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�l�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����P��N1�����
�b�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�g�<�3��e�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
�9�
�0�8��(�������l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�o�(���@�ӓ�F��d:��9�������w�m��������l�N�����u�8�f�
�"�d�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�g�
� �n�m����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���3�
�g�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��M���
�f�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�CU��Q��@؊�g�o�����4���:����V��X����n�u�u�&�0�<�W�������D9��hW�*��o������!���6�����Y��E��u�u�&�2�6�}�(�������T��^1��*���
�g�o����0���/����aF�
�����e�n�u�u�$�:��������_	��Y�����c�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����l��X�����;�!�3�
�`��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��U�����<�<�;�!�1��Aׁ�K����g"��x)��*�����}�u�8�3���B�����Y�����`�
� �l�d�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E����� �l�e�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���d�e�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G]�����e�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӗ��R
��1�����
�m�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������V
��Z�*���l�m�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƹ�l��x��Gӊ�:�4�
�
�"�l�Fف�J����g"��x)��*�����}�d�3�*����P���F��P ��U���-� �,� ��(��������U��\�����u��
����2���+������Y��E��u�u�&�2�6�}��������l*��G1�*ڊ�
�
� �d�e��C��*����|!��h8��!���}�e�1�"�#�}�^�ԜY�ƿ�T����*����'��:��d�G���I�ԓ�F9��W��D��������4���Y����W	��C��\�ߊu�u�<�;�;�<����&����	��h_��G���e�3�
�e�n�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�f��(���&����lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���?����\	��W��*���
� �d�a��o�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�����'��:�
�n�o����K����V��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�6�/��������\��1�����a�3�
�d�b�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����g�
�0�o���;���:���F��P ��U���'�!�'�
��/���*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��^	��ʴ�
�0� �;�f�-����Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�D�����%�'�!�'������Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������4�
�0� �9�n����Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����u�%�'�!�%��(�������g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����9�4�
�0�"�3�B�������`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����4�u�%���.�W���-����t/��a+��:���`�1�"�!�w�t�}���YӅ��C	��Y��3җ�d��3�e�1�(�(���
����@9��h_�����&�u��u�w�:������ƹF�N��1������]�}�W���Y����`2��rN�<�����_�u�w�}�W���I����g.�'��0���n�u�u�u�w�9�ށ�0����	F��c+��'�ߊu�u�u�u�8�)� ���1����}2��r<��N���u�%�'�u�]�}�W���Y����\��yN��1��������}�D�������V�=N��U���u�<�d�o��}�#���6����e#��x<��F���:�;�:�e�l�}�W���Yӂ��GF��x;��&���������W��Y����G	�N����u�;�u�:�'�3���s�����G�������d��1�m��������]��1�<�ߊu�u�0�0�>�}�}���Y���z"�'��0���n�u�u�u�w��:���8���/��r)��N���u�u�u�1�9��>���Y�ƅ�g#��eUךU���u�u�:�!� ��?��0����v4�d��Uʥ�'�u�_�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u�%�.���0�Ɵ�w9��p'�����u�u�u�<�g�g�>���-����t/��a+��:���c�u�:�;�8�m�L���Y�����N��U���
���n�w�}�W�������	F��cN��1��������}�D�������V�UךU���;�u�:�%�9�3�L�ԶY����\��Y��U����d��3�g�;����J����R��'��U���2�;�'�6��}�W���Yӯ��	F��c+��'�ߊu�u�u�u���#���Y�ƅ�g#��eUךU���u�u�<�e� ��?��0����v4��N��U���1� �
���}�W���<����]ǻN�����}�u�u�u�w�9����Y����g"��x)��*�����}�d�3�*����P���F�N�� ���u� �u����>���<����N��
�����e�u�n�u�w�8�Ͻ�����]��=d�����_�u�u�
��0�������]��1�����1�%� �u�w�2�����ơ�$��*��*ڊ�8�9�f�;��o���&¹��K9��Gd��Uʲ�;�'�6�8�'�u�W���Y����wF�_�U���u�u�����2��Y��ƹF�N��������h�w�o�}���Y���W��h9��!���k�f�y�u�w�}�WϺ�����w2��
P��G�ߊu�u�:�!�:�-�_���Y�����N��U���-� ���#�o�(���K�ޓ�JǻN��U���<�d�h�u��%�"���6���� 9��h\�*��_�u�u�u�w�2���Y����~3��N!��*���3�
�d�
�e�f�}���Y����@��Q��A���f�
�
�d�w�}��������^ ��_��A���
�<�:�%�a�3�(���K�����R��U���u�_�u�u�w�}�3��Y��ƹF�N�� �����u�k�e�W�W���Y�ƨ�]V��~*��U��c�y�u�u�w�}����&����{F�]����u�:�!�8�'�u�W���Y����_�	N��*���y�u�u�u�w�/����D�ƭ�l��d��U���u�1�;�u�i�:����&����CV�N��U���6�u�k�2�'�;�(��&����F�N�����u�k�2�%�1��E݁�H��ƓF�Q1�����!�f�;�
�c�l�"��CӅ��C	��Y��3җ�d��3�e�1�8�������lWǻN�����<�u�4�u�]�}�W���Y���F��=N��U���u� �
���}�I��s���F�S��*����u�k�f�{�}�W���Yӂ��G9��s:��H���a�_�u�u�8�)����Q���F�
��E��u�
�&�<�9�;�(��&����F�N�����u�k�1�4�$�:�(���K�ӓ�O��=dװ���u�x�!�0�4�/����
����N��h-�����u�3�!�0�$�<�ϳ�����F�=N��U����
�&�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���	����U��S�����
�!�
�&��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����s���F�N��U���u�u�4�
��;���Y����`9��ZUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W������G��h^�����4�&�2�u�%�>���T���F��h�� ���e�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���	����F��1�����h�4�
�:�$�����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C]�����|�4�1�;�#�u��������F9��1��U���%�6�;�!�;�l�G���PӒ��]FǻN��U���u�u�u�u�w�}��������9��R	��Hʴ�'�9�
�:��2���&����9��E��D��_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����E�����
�'�2�4�$�:�W�������K��N�����0� �;�d�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���R��R�����%�0�u�h�6�����&����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9����Q����P	��h��G���%�u�u�%�4�3����H���O��_�����u�u�u�u�w�}�W���Y����V��Y1�����u�h�4�'�;���������
9��R1�����d�e�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F������'�
�
�'�0�<����Y����V��C�U���4�
�0� �9�o����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�V�����;�g�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�������V��T��*���g�a�%�u�w�-��������lV�G�����_�u�u�u�w�}�W���Y���R��R�����%�0�u�h�4��9���8����A��1��E���2�d�c�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C�����!�'�
�
�%�:�����Ƽ�\��D@��X���u�4�
�0�"�3�D�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��*��� �;�f�%�2�}�JϿ�&����G9��\��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ�ӈ��N��^����� �g�a�%�w�}��������EW��G��U���;�_�u�u�w�}�W���Y���F��h�� ���f�%�0�u�j�>�(���<����G��hZ�����'�2�d�g�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���'�!�'�
��/�Ͽ�
����C��R��U���u�u�4�
�2�(����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N�����0� �;�a�'�8�W������]��[�*��u�u�u�u�w�}����s���F�N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!��.�(�������\�R�����
� �g�a�'�}�W�������l
��h^��\���=�;�_�u�w�}�W���Y���F�V�����;�a�%�0�w�`����7����a4��E��C���e�'�2�d�c�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���%�'�!�'����������]F��X�����x�u�u�4��8����L����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʴ�
�0� �;�b�-����DӇ��P	��C1��F؊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�����PӇ����F�����;�
� �g�c�-�W���	����@��A_��\���u�=�;�_�w�}�W���Y���F�N��*��� �;�`�%�2�}�JϽ�&����k'��C��*���0�d�'�2�f�i�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u��9�
�8�����
����lT�������%�:�0�&�w�p�W�������l ��h"�����'�2�g�c�6�.���������T��U´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������W������u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���u�u�u�u�>���������C9��E��G��i�u��9��2�(���	����A��_�N���u�u�u�u�w�}�Wϻ�
�����T�����2�6�d�h�6�����
����g9��1����|�!�0�u�w�}�W���Y���F�N��9���
�:�
�:�'�.����K���F��h�����#�
�n�u�w�}�W���Y����������u�u�u�u�w�3�W���Y���F���U���_�u�u�;�w�/����B���F������%�:�0�&�w�p�W���	����@�V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���H����[��N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�(���&�����Yd��U���u�u�u�u�w��(���&����Z�q\�� ��m�%�n�u�w�}�W���Y�����GY�����g�l�i�u�4�-�(���J�֓�]ǻN��U���u�u�u�u�$�8�(���&����Z�^��*��� �f�m�%��n��������]ǻN��U���u�u�u�u�:��N�������F���*���3�
�a�
�e�W�W���Y���F�N����
�0�
�g�e�a�W���&�ԓ�F9��1��N���u�u�u�u�w�}�WϪ�	����A��_�U��!�%�`�
�"�n�O���B���F�N��U���u�8�
�e�%�:�F��Y����^��1��*��
�f�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=N��U���4�&�2�u�%�>���T���F��X�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������A��N���ߊu�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�ӓ�@��G�����_�u�u�u�w�}�W���Y����VW��[�����g�<�d�
�2��E��E�ƞ�]��h��*���&�g�<�d��(�N���	��ƹF�N��U���u�u�0�0�2�����&����T��R�����!�1�/�'�$�;�(��&����F�N��U���u�u�;�"�>�3�������� S�
N��#���
�
� �c�a�-�_������\F��UךU���u�u�u�u�w�}�(���K�ӓ�V��\�I���
�4�g�`�1��Aف�J���F�N��U���u�!�%�f��8�(��I���G��W�� ��c�%�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�&�<�;�'�2����Y��ƹF��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G��U���;�u�u�u�w�}�W���YӇ��l
��q��9���
�l�g�0�g�k����H���F��E1��*���
�:�%�d���(߁�&����Q��G]�U���u�u�u�u�w�}��������A9��X��L���0�d�'�2�f�m�K�������l ��h"����
�
�
�
��(�F��&����F�N��U���u�u�6�
���6�������9��1����c�i�u�'��)�1���5����_��h��*ي� �d�b�
�d�W�W���Y���F�N��*������0�:�i�(���&����^��S�����!��'��8��N����ד�l ��^�*��_�u�u�u�w�}�W���Y����}"��v<�����a�
�
�
�2��D���DӇ��l
��q��9���
�l�g�0�g�l����I�Г� ]ǻN��U���u�u�u�u�;��3���+����^9��h��*���
�l�u�h�6�/��������\��1�����`�3�
�d�e�-�L���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�u�u�x�w�.����	����@�CךU���'�6�&�u�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H��r�u�=�;�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�����d�|�u�=�9�}�W���Y���F������
�0�8�l��8�(��M���T��Q��G؊�d�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǻN��Xʴ�&�2�u�'�4�.�Y��s���C��R��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������A�C�����u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���J����lT�V ��]���!�:�1�3��n�(��DӇ��P	��C1��D��|�u�=�;�w�}�W���Y���F��d1�� ����!�g�
�2��F��E�ƪ�l��{:�� ���f�3�
�d��o�}���Y���F�N�����!�%�
�0��l�B��Y����G��h��G���%�n�u�u�w�}�W���Y����V
��Z�����d�b�i�u�2���������l��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}���Y���R��P �����&�{�x�_�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�f�1�0�E���Y����9F�N��U���u�u�u��;���������9��P1�@���h�<�
�<��/�;���&�ד�F9��1��N���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B���F���U���!�&�4�0��-�9���
����UF��RN�����8�6�<�0�w�p�W�������l ��h�����%�:�u�u�%�>��������R����6���&�y�4�
�2�}��������F9��1��\���u�7�2�;�w�}�W�������R��d1��ʼ�_�u�u�u�w�}�W���Ӈ��`2��C_�����u�k�_�u�w�}�W���Y���Z �F��*���&�
�:�<��}�W�������]��X�����!�'�u�u�'�>��������lV�G�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�e�;���s���F�N��U���0�&�_�u�w�}�W���Y���F�V��&���8�i�u�%���ށ�
����9F�N��U���u�u�u�;�w�;�}���Y���F�@��U����
�!�
�$��W���s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�D�������F�N��U���u�u�0�&�]�}�W���Y���F�N������3�8�i�w�-�$�������^9��=N��U���u�u�u�u�w�3�W���s���F�N�����u�%��
�#�����Y���F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u��������U��Z��G��4�
�:�&��+�(���P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y���F��[��U���4�
�:�&��2����Y�ƭ�l����U°�<�6�;�
�"�o�C���Y�ƭ�l��D��ۊ�|�|�!�0�]�}�W���Y���F�N������3�8�i�w�-�$���ǹ��^9��=N��U���u�u�u�u�w�1����Y���F�N��U���u�%��
�$�}�JϿ�&����GU��D��N���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�=�;�4��	��������[�=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���4�
��3�:�a�W���*����9��Z1����u�u�u�u�w�}�W������F�N��U���u�u�u�%������DӇ��`2��CZ�����n�u�u�u�w�}�W���YӃ����=N��U���u�u�u�=�9�<�(���
�ӓ�@��S����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�4�
��;���Y����g9��1�����_�u�u�u�w�}�W���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:��ߊ�&�
�n�u�w�}�W���Y����������u�u�u�u�w�5�Ͽ�&����GP��D��U��_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�6��$������R��c1��F���8�g�_�u�w�}�W���Y���V
��=N��U���u�u�u�u�w�}�W���7����^F���&���!�
�&�
�l�}�W���Y���F���U���_�u�u�u�w�}�W���Ӊ��V��
P�����u�u�u�u�w�}�W���7����^F�L��-���w�_�u�u�w�}��������F�R �����0�&�_�u�w�}�W���K����G9��hZ�*��i�u�!�
�8�4�(�������V��RF�����}�g�g�3��i�(��U���lǻN��G���3�
�a�
�d�a�W���Y��� ��E��D��u�=�;�}�:��G���&����CT�N��R��u�9�0�_�w�}�W�������l ��]����u�u��
�"�n�O���Y����G��X	��*���!�'� �&�0�8�_�������l
��1�F���u�;�<�;�3�)��������9��G�U����;�0�
�;�����H����R��G\��H���8�f�
� �`�m�����Ƹ�C9��h��B���%�|�_�u�w�<��������]��1��DҊ� �l�a�%�w�`�_�������Z9��hX�*��4�1��;�2���������l��B1�G���|�_�u�u�6�:�F�������@9��^1��*��
�f�i�u�w�}�W���+����9��[1����� �m�a�%�w�5��������W_��^1��*��
�g�e�u�w�l�^ϻ�
��ƹF�N�����8�g�
� �o�i���Y����R��1�����0�
� �m�c�-�W��Q����VT��[�����d�<�3�
�g��DϿ�Ӵ��T��V�����
�
� �b�a�-�^�ԜY�ƞ�]��h��*���:�
�
� �o�i����D������YN�����
� �a�f�'�}�W�������l
��1�U���0�w�w�_�w�}����H����l��X��*��� �m�m�%�w�`�}���Y���C9��h�� ��g�%�u�=�9�u��������Z9��hV�*��e�u�u�d�~�8����Y���F��R����
� �m�e�'�f�W���+����9��[1�����3�
�g�
�e�a�Wǌ�����R
��X ��*ۊ� �b�c�%�w�2�W�������l
��h_����u�4�2�g��l����A����Z�D�����6�#�6�:��5��������F��P ��]���
�
� �a�d�-�^ê�&����T��B �����}�e�u�u�:��B���&����CW�C����!�u�|�|�~�W�W�������l��h�����<�3�
�e��n�K���Y���F��V ��G���9�:�0�
�"�j�C���Y����N��h�����<�3�
�b��o�G���Y�����RNךU���u�u�0�d�1��A߁�K���F��Y	��*���
�;�&�3��d�(��E���F��R ��'���0�
�
�
�"�j�E���Y�ƾ�e9��hY�*��u�9�0�w�u�W�W���T�ƭ�l��RN�����u�'�6�&�y�p�}���Y����\��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����VJ��G1�����0�
��&�d�;���Y����P	��h��G���%�|�u�u�5�:����Y�����F�����4�
�:�&��2����Y�ƭ�l��E��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^�������C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*���� 9��Z1�U���u�:�}�0�>�>��������l��
N��*���&�
�#�
�~�t�^Ϫ���ƹF�N��U���%�1�;�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��X ��I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���0�4�&�2�w�/����W���F�V�����4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�N�����;�u�u�u�w�4�W�������C9��Y�����6�d�h�4��)����Y������T�����2�6�d�h�6�����
����g9��1����|�u�=�;�]�}�W���Y���R��S��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�<�(������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������R��V�����'�6�&�{�z�W�W���	����W��D�����:�u�u�'�4�.�_�������C9��P1������&�f�3�:�o�W�������l ��]�����u�u�7�2�9�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1����u�;�u�:��8��������lT��h�Hʴ�
�:�&�
�!��^���Y����l�N��U���u�4�
�0�3�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���%�'�!�'��}����Ӗ��P��N����u�%�'�!�%��(�������A	��N�����&�4�
�0�w�-��������`2��C]�����y�0�<�6�9����M������h��3����:�
�l�e�8�G�������^�V�����;�e�%�0�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�f�3�8�e�}��������K��X �����f�
�g�h�6�����&����O�N�����u�u�u�u�w�}��������lV�
N�����
�:�
�:�'�l�(݁�&ù��A��[����u�u�u�9�2�W�W���Y���F��h�� ���e�i�u�%�%�)����&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�0� �9�l�����Ƽ�\��D@��X���u�4�
�0�"�3�F���
����C��T�����&�}�%�6�{�<�(���&����l5��D�����g�u�-�!�8�9����Jǹ��F��E1��*���
�:�%�d���(ށ�����J��G1�����
�
�'�2�]�}�W������F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<�ϰ��Ω�Z��Y
�� ��a�%�u�u�'�>�����ד�O����ߊu�u�u�u�w�}��������F���*����'��:��d�E���H����lW��d��U���u�0�&�u�w�}�W���Y����C9��C��*���h�4�
�0�"�3�F�����ƹF�N�����3�u�u�u�2�9��������9l�N�U���'�!�'�
�w�.����	����@�CךU���%�'�!�'����������PF��G�����4�
�0�u�'�.��������l��h��*���0�<�6�;��(�E���	����_9��s+��'���'�
�a�0�g�/���O�ƭ�l��B��G���0�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��F���8�g�u�;�w�2�_ǻ�����W9��h\�*��h�4�
�:�$��ށ�P���G��d��U���u�u�u�4��8����K���P
��y*��4���0�8�a�
������M��ƹF�N�����_�u�u�u�w�}�W�������]9��S�����!�'�
�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h�� ���f�4�&�2�w�/����W���F�V�����;�f�4�&�0�����CӖ��P�������4�
�<�
�$�,�$�������^9�������1�3�
�f��o�W���0����r4��R��Aފ�
�
�0�
�o�q��������lU��E�����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GU��D��\ʴ�1�;�!�}�/�)��������9��S�����;�!�9�d�g�t�^Ϫ���ƹF�N��U���%�'�!�'��}�JϽ�&����k'��C��*���0�d�'�2�f�o�}���Y���V
��d��U���u�u�u�4��8����J���R��R�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������G��hZ�����;�%�:�0�$�}�Z���YӇ��A��E ��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�n����K�Ʃ�Z��Y
�� ��a�%�y�6���2���+����lR��R1�����d�a�u�%�%�)����&����l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����0�<�6�;��(�E���	���R��X ��*���
�|�|�u�?�3�}���Y���F�V�����;�a�i�u�;��3���+����^9��h��*���
�f�n�u�w�}�Wϻ�
��ƹF�N��U���%�'�!�'��}�JϿ�&����A��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������R��P �����&�{�x�_�w�}��������9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�
�&��q��������U��Z��G���9�����)����O����l��h_�Yʴ�
�0� �;�b�-����Y����V��=N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�d�;���Y����]	�������1�3�
�f��o�JϿ�&����G9��1�\���!�0�u�u�w�}�W���YӇ��A��E ��U��6�
��������MŹ��9��P1�A�ߊu�u�u�u�;�8�}���Y���F�V�����;�`�i�u�'�/����&ƹ��V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h_�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�a�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h_�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�`�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(������]F��X�����x�u�u�4��4�(���&�ғ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��N�U´�
��3�8�g�9� ���Y�����T�����d�d�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�h�W�������A	��D�X�ߊu�u�%�&�0�?���&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����^�
N�����;�!�9�d�f�`����*����W��X����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�c�<����Y����V��C�U���4�
�<�
�3��C���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������[�V�����
�#�
�u�w�-�4���
����W	��C��\��u�u�0�1�'�2����s���F������7�1�l�u�$�4�Ϯ�����F�=N��U���&�2�7�1�n���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����M�����T�����d�d�h�4������Jӂ��]��G����u�;�u�'�4�.�L�ԶY���F��h��*���$��
�!��.�(���
������T��[���_�u�u�%�$�:����&����GW��D��*���<�;�%�:�w�}����
�έ�l��h��*��_�u�u�0�>�W�W���Y�ƥ�N��h��*���
�a�u�=�9�W�W���Y���F��h��*���$��
�!��.�(���DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����<�
�&�$���ށ�
����[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�ƭ�l��h�����
�!�
�&��}����Ӗ��P��N����u�%�&�2�4�8�(���
�ԓ�@��h�����%�:�u�u�%�>����	����l��h[����u�0�<�_�w�}�W����έ�l��h��*��u�=�;�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��F1��*���
�&�
�u�$�4�Ϯ�����F�=N��U���&�2�6�0��	��������l��^	�����u�u�'�6�$�u��������lQ��=N��U���<�_�u�u�w�}����	����l��hY�U���;�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������B9��h��*���
�u�&�<�9�-����
���9F������6�0�
��$�i����J����Z��G��U���'�6�&�}�'�.��������9F����ߊu�u�u�u�1�u��������l_�����ߊu�u�u�u�w�}��������B9��h��*���
�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����Z��D��&���!�
�&�
�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�.��������l��h��*���&�<�;�%�8�8����T�����D�����
��&�`�1�0�C���
����C��T�����&�}�%�&�0�?���O���F��P��U���u�u�<�u�6���������O��_�����u�u�u�u�w�-��������`2��C[�����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GP��D��U���<�;�%�:�2�.�W��Y����C9��P1������&�c�3�:�h��������\������}�%�&�2�5�9�F��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��h��*���h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���
����@��d:��܊�&�
�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���'�
�!��%�����@�֓�lV��h��D��
�d�i�u�#�����&����\��R�� �&�2�0�}�%���������C9��h^��*ڊ� �d�g�
�c�q�E���s���R��[�����:�%�d�
���(���H����CR�
N��*�����!��5�/����O����V��h�F���:�;�:�d�l�}�WϿ�����u	��{��*���e�0�d�3��m�D���Y����G��X	��*���!�'� �&�0�8�_���&����\��X��Dӊ�
�
�
�
�"�l�Dց�H���F��P ��]��� �g� �
�n�1����/����V��h�\�ߊu�u�'�
�#���������lT��h^��*���d�`�
�f�k�}�W���Y����_9��s+��'���'�
�c�0�g�/���Mӑ��]F��R�����'�2�d�c��t�J���^�Ʃ�@�N��U���4�'�9�
�8�����Hʹ��V9��Q��E���%�n�u�u�6�/��������\��1�����g�3�
�e�d�-�W��s���F�V�����:�
�:�%�f��(���&����lW��1��U���;�}�0�
�:�����H���F�_��U���0�_�u�u�w�}����=����a��Z1�*���
�0�
�a�l�}�WϿ�����u	��{��*���g�0�e�f�1��G���	���l�N��Uʶ�
�����8���&����A��Z����u�&�9�!�'�����H���F�_��U���0�_�u�u�w�}��������l*��G1�*؊�
�
�
� �f�k�(��s���R��[�����:�%�d�
���(ځ�����9��R�����u�u�u�'��)�1���5����_��h��*؊� �d�f�
�f�*����
����^��E��D��}�|�h�r�p�}����s���F�V�����:�
�:�%�f��(���&Ź��T9��UךU���'�
�!��%�����@�ԓ�lV��B1�Aӊ�f�i�u�u�w�}�WϽ�&����k'��C��*���0�e�'�2�f�i� ���Yە��l��h��*��b�e�u�u�f�t����Y���F���*����'��:��d�G���I�ԓ�F9��W��D�ߊu�u�'�
�#���������lT��h_��*���d�m�
�f�k�}�W���Y����A��C1�����:�
�l�e�2�l����I�Փ�F��R �����!�%�
�0��l�B��Y���O��[�����u�u�u�'��)�1���5����_��h��*���
�b�n�u�w�<����&����	��h_��G���d�g�3�
�g�l����D���F�N�����
�:�
�:�'�l�(߁�&¹��lW��1��U���;�}�0�
�:�����H���F�_��U���0�_�u�u�w�}����=����a��Z1�*���
�0�
�m�l�}�WϿ�����u	��{��*���g�0�d�f�1��G���	���l�N��Uʶ�
�����8���&����A��V����u�&�9�!�'�����H���F�_��U���0�_�u�u�w�}��������l*��G1�*؊�
�
�
� �f�d�(��s���R��[�����:�%�d�
���(ہ�����9��R�����u�u�u�9���/�������P��h_�����l�u�=�;��8�(���&����W��^��H��r�u�9�0�]�}�W���Y����_��X�����d�
�
�
��(�F��&����F�V�����:�
�:�%�f��(���&ƹ��lW��1��U��_�u�u�u�w�1�>���!����V��X��*ۊ�0�
�l�u�?�3�_���&����l��h_�@��u�u�d�|�2�.�W���Y�����h��3����:�
�l�e�8�F�������S��UךU���'�0�2�
�"�d�G���Y���F��E�����!�3�
�c��o����&�ѓ�V��P�����!�3�
�b��o�L���Yӄ��V��h��*���
� �l�m�'�}�J���&�ѓ�V��P�����
�`�
�g�6�9��������l��h��L���%�|�_�u�w�<����&����lP��h�I���&�9�!�%�g�;�(��&����]��Z��M���
�g�
�g�l�}�WϺ�����]9��h\�*��i�u��-��	�8���K����T9�� [�U���1�9�!�1�-�/����&����CU�
NךU���u�u�4�2�f�<��������Z9��hV�*��"�0�u�6�%�$�F�������9��^��H��r�u�9�0�]�}�W���Y����VW��[�����
�
�
� �o�e���Y����K��X �����f�
�g�i�w�l�W����Υ�l
��q��9���
�
�0�
�g�}�W�������l
��h]�����u�e�n�u�w�8����	����F9��1��U��<�0�
�
�"�n�O���Q����\��XN�\�ߊu�u��-��	�8���K����lT��h�I����;�1�
�2�0�N߁�����R��N�������,� ��n����H˹��Z�=N��U���u�;� �0�4�3�(������@��C��*���g�m�%�}�~�`�P���Y����l�N��Uʦ�9�!�%�
�"�o�E���B���F�	��*���g�g�6�u�$�4�Ϯ�����F�=N��U���
� �g�g�4���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�%�6�{�<�(���&����l5��D�����d�_�u�u�2�4�}���Y���Z �F��*���&�
�:�<��}�W�������]�F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�3����	����A������!�9�2�6�g�t�W���Q����\��h�����u�u�%�&�0�>����-����l ��h_��\���=�;�_�u�w�}�W���Y����U��\����u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}��������9��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��ԶY����A��B1�G���u�h�&�1�;�:��������A��M�����;�1�<�
�2�4���U���l�N��*����'��:��l����Mù��Z�D�����6�#�6�:��3����ۏ��_��X�����&�'�2�g�a�}�W���������T�����g�d�|�_�w�}����&����V��N�U��u�=�;�}�>�3�Ǫ�	����U��^��A���u�<�;�1�6�����&����lV������w�_�u�u�4�-����N¹��Z�_�����u�!�%�`��(�C���	���R��X ��*���
�|�0�&�w�m�L���Yӏ��T9��Q��EҊ�d�i�u�
�$�4����&����CW��N����� �b�c�%�w�`����M����lQ��h�D���d�1�"�!�w�t�}���Y����e9��Q��D݊�g�i�u�!��2����������^	��´�
�:�&�
�!�i�G���Y����T�������!�d�
� �c�n����B�����h8�� ��f�%�u�h�]�}�W���Y����e9��Q��D݊�g�"�0�u�>�3��������N��S��D���0�&�u�u�w�}�WϮ�+����G9��h��A���%�n�u�u�8�����H����F9��1��U��}�8�
�a�1��Aف�KӇ����1��*��
�g�n�u�w�2�(����Փ�l ��^�����h�}�8�
�c�;�(��&����]��R�� ��e�%�|�_�w�}�(�������S��G\��H���4�2�d�4�;�'����H����R��G\��ʧ�#�3�
�g��o�L���YӖ��9��Z�����
� �l�b�'�}�J�������U��\��Gʺ�u�0�0�0��8��������P�=N��U���b�1�8�'�6��(���&����R��N�U¥�l�
�0�:�0�3����&����CT��X�����;�!�9�d�f�f�W���	����Z9��hV�*��i�u�!�%�c����I����R��e��ۊ�9�
�0�:��(�O���	����F�G1�����
�f�3�
�f��F��Y����_	��T1�����}�0�<�0�"�.����Q����^��B1�C���|�`�|�n�w�}����
����@9��h[�*��i�u�8�;��;�(��&����]��Z��F���
�`�
�g�l�}�WϮ�/���� 9��h[�*��i�u�u�u�w�}����LŹ��lS��h����u�!�%�g��(�C���	����[�I�����u�u�u�u�w�.��������U��[��F�ߊu�u�
�4�e�i����Iʹ��Z�D�����6�#�6�:��3����ۖ��R
��1��*��
�f�u�u�9�4��������9��hX�*��|�_�u�u��<�E�������9��R�����u�u�u�0��0�Fށ�����l��@��U¦�9�!�%�a�3�0����&����W��F�U���d�|�0�&�w�}�W���Yӕ��A��E	�����
�m�
�f�]�}�W����ԓ�l��h��L���%�u�h�_�w�}�W���&����lS��R	��G��"�0�u�7�:�/��������l ��X�����|�h�r�r�w�1��ԜY���F��h�����#�g�����L���YӖ��C9��h]�*��i�u�!�
�8�4�(�������]��Y�����`�
� �f�o�-�^�������]��V�����
�#�
�|�l�}�W���YӖ��9��D�� ��`�%�u�h�$�9��������G	��E�����<�;�1�%�$����I����U��UװU���%�&�
� �a�m����Dӕ��l
��^�����'� �&�2�2�u�E�������O������1�4�
�:�$�����K���9F�N��U���g�6�&�
�"�k�C���Y����G��X	��*���!�'�'�&�-�u����ۖ��9��hX�*��y�g�|�_�w�}����&����_��N�U���
�:�<�
�2�)�ǫ�
����WN��h��*��d�u�u�;�>�3�ǿ�&����G9��\��D���_�u�u�7�6�.����&����
_��N�U§�<�<�3�
�n��EϿ�ӗ��U��\��F��u�u�$�
�"�h�E���Y���F�N�����2�'�2�d�o�}����Q���� V��B1�E���}�|�h�r�p�}����s���F�C��@݊� �`�a�%�l�}�WϬ�/����^��G\��Hʦ�1�9�2�6�!�>��������A��CF�����0�}�%�6�9�)���&����u ��q(��3���!�
�;�0�2�u�������A���*���3�
�b�
�f�n�Z�������V�G����u�
� �`�a�-�W��Q����9��P1�D���;�u�8�
�a�;�(��&���9F���*��� �`�f�%�w�`�_���&�Г�F9��1��U���'�3�
�b��o�L���YӔ��9��hY�*��i�u�!�%�`����K����K	��V�����
�#�
�|�]�}�W���&����V��N�U¡�%�c�
� �`�o�����ƭ�l��D��ۊ�|�_�u�u�2����&����Q��N�U¡�%�3�
�a��o��������9��hZ�*��n�u�u�&�;�)�������� 9��R�����u�u�u�
�6�o�C���&����CT��_��]���
�8�d�
�"�k�@���Q���A��N�����u�u�u�u�$�1����&����_��UךU���0�
�8�d��8��������P��G\��H���8�
�g�'�0�l�F���Ӓ��lT��Q��Fڊ�g�n�u�u�$�1����&����T��N�U���u�u�u�<��-��������[����*���
� �g�c�'�u�^��^���V
��d��U���u�<�
�%�%�8���s���@��C��F���
�c�
�g�k�}����Oʹ��lQ��h����8�
�a�;�#�;�(��&���9F���*���g�
� �m�o�-�W��Q����^��B1�M���u�;�u�0��0�E܁�����l��d��Uʦ�9�!�%�`�1��@ہ�J���9F�N��U���2�d�4�9�8�8�(ށ�����l��@��U¦�9�!�%�a�1��Aׁ�K���F�G�����_�u�u�u�w�8�(���N�֓�]ǻN�����8�g�
� �o�m����D���F�N�����
�9�
�0�8����O����D��F�����%�a�3�
�a��E��Y���O��[�����u�u�u�
�b�4����Lù��l�N�����%�b�3�
�e��E��Yے��lU��E��D��u�:�u�%�4�3����H���9F���*���g�
� �l�b�-�W��Q���� 9��hW�*��4�1�<�;�0�/���A����F�D�����l�3�
�a��o�K�������
9��P1�A���;�u�&�0��8�(��I��ƹF��R�����3�
�`�
�e�a�W��Y����N��h��3����:�
�
�2��G���Y����\��h��*���0�&�u�e�l�}�Wϭ����� V��B1�M���u�h�_�u�w�}�W�������l
��1����u�!�%�`��(�N���	����[�I�����u�u�u�u�w�-�!���&ƹ��T9��W�U���&�9�!�%�f�;�(��L����[�C��Dӊ�0�
�d�`�/�/��������_��G�U���&�9�!�%�e�;�(��I����[�U�����3�
�m�
�e�<�ϭ����� W��B1�Eߊ�g�n�u�u�$�1����&����_��N�U���u�u�u�!�'�h�(���M�ד�F��R �����g�
�0�
�e�o�G���Y�����RNךU���u�u�
�4�e�i����Iʹ��l�N�����%�
� �c�a�-�W��Q����T��R	��G��-�'�4�
�8�.�(���&����F�D�����3�
�a�
�e�a�W��Y����N��h��3����:�
�
�2��G���Y����\��h��*���0�&�u�e�l�}�Wϭ�����A��Q��Eߊ�f�i�u�u�w�}�WϿ�&����G9��\��3�����"�0�w�4��������^��G��U��|�0�&�u�w�}�W�������]��[�*��u�u�&�:�2�8����&����U��N�U���u�u�u�!�'�o�(���M�ѓ�F��R �����
� �a�d�'�u�^��^���V
��d��U���u�4�
�:�$�����I���F��G]�����a�
�g�i�w�1�(���N�Г�F��SN�����
�g�
�g�l�}�WϪ�	�Փ�F9��1��U��}�0�&�2�5�)����H����R��D�����b�3�
�g��o�L���YӒ�� R��B1�G���u�h�}�&�2�����H����AF��[1�����3�
�g�
�e�f�W�������9��hZ�*��i�u�4�
�8�.�(���&���G��]�����d�e�n�u�w�)���&����T��N�U��u�=�;�}�:��@���&����CW������!�9�c�
�~�8����I��ƹF��Z��E���
�f�
�g�k�}�F������@��R
��G���2�d�e�|�i�.����Q����\��h��G��|�0�&�u�g�f�W�������9��hZ�*��i�u�!�
�8�4�(�������]��Y�����:�&�
�#�e�m�W�������V��1����e�|�n�u�w�)���&����R��N�U��u�=�;�}�/�����&����R��N�����:�&�
�#�f�i�D������D��N�����g�
� �a�b�-�W��[����[�������1��
�
�"�i�G���P����]��Y�����:�&�
�#�e�n�^������D��N�����g�
� �a�`�-�W��
����\��h�����&�<�!�9�1�u��������^��1��*���
�d�y�:�>�)��������]��^��Sʓ�
�
�4�!�1��C؁�H����F��@ ��U���|�|�_�u�w�0�(�������9��R�����9�2�6�#�4�2�_�������]��Y��3؊�
�4�!�3��i�(��U���l�N����
� �a�`�'�}�Jϭ�����Z��R��¦�<�!�'�2�#�.����Q����e9��hZ�*��y�:�<�!�0�/��������V�N����
� �a�d�'�u�F������\F��G��N���u�!�%�f��(�B���	���D�������<�;�1���8�(��H���@��R
�����;�!�9�d��k�^ϻ�
���]ǻN�����d�3�
�g��o�K�������T��A�����;�<�;�1������K���F��D�����%�6�;�!�;�l�(���P��ƹF��Z��F���
�b�
�g�k�}��������E��X�����;�1��
�"�n�O���P����]��Y�����:�&�
�#�e��2���s���G��Z�� ��g�%�u�h�u�� ���Yە��]��C��Fي� �f�c�%�~�c�����έ�l��D�����f�|�u�9�2��U�ԜY�Ƹ�C9��h��@���%�u�h�w�u�*����	����F
��D1��*��
�g�h�4��2�����ғ�F��D��D��u�u�!�%�d����L����[��C
�����
�0�!�'�%�.��������V��U1�����
�
� �`�n�-�^��P��ƹF��Z��M���
�g�
�g�k�}����OĹ��lP��h����4�
�:�&��+�(���s���G��W�� ��c�%�u�h�u�� ���Yە��]��G��*���c�e�%�|�k�.����Q����\��h��G��|�u�9�0�u��}���Y���G��_�����3�
�f�
�f�a�W���&����P9��T��]���<�0�&�2�2�u����H����T��G\��F���n�_�u�u�:��F���&����CW�
N�����2�6�#�6�8�u����ۓ��Z��SF��ۊ�4�!�3�
�o��F��M����F�C��A؊� �b�e�%�w�`��������l��C�����!�'�2�!�$�:��������U��]��F���:�<�!�2�%�(�������F�C��Aۊ� �b�c�%��l�FϺ�����O�G�U���!�%�a�
�"�j�A���Y���D��_��]���;�1�%�&��(�A���	�����Y�����:�&�
�#�e�n�^������D��N�����a�
�:�
�"�e�A���Y���G��Z�� ��c�%�u�:�w�-��������lW�=N��U���
�`�3�
�`��F��Y����_	��T1�����}�0�<�0�"�.����Q����l��C1��*��
�d�y�a�~�W�W�������l ��\�����h�w�w�"�2�}�%�������9��hY�*��h�4�
�:�$�����I�Ʃ�@�L�U���!�%�a�
�"�n�E���Y����A��a1��*��
�d�c�u�w�}�������9F���*���3�
�f�
�e�a�W��Y����N��D\�� ��l�%�u�u�'�>�������� P�R��U��n�u�u�!�'�i�(���@�֓�F�F�����
�9�
�;�$�o���&����T����U���6�;�!�9�f�l�L���YӒ��lS��Q��Lي�g�i�u�!�'�l�(���&����	��B �����"�3�
�a��n�L���YӒ��lS��Q��FҊ�d�i�u�'�0�����I˹��S��N����!�u�|�_�w�}����M����S��G_��Hʸ�;��3�
�e��D��Y����W	��C��\�ߊu�u�8�
�b�;�(��&���F��h\�� ��e�%�}�d�3�*����P���F��G1�*���`�d�%�u�j�)���&����
S��F�U���u�:�;�:�g�f�W�������9��h[�*��i�u�4�
��(�C���	�θ�l��R	��]���<�;�1�!�'�i�(�������U��G_��U���;�:�!�
�9�8��������V��Z��D���&�
� �`�g�-�^���������^ ����� �&�2�0��0�(�������U��^��D���h�e�4�1�#������ι�@��R
�����d�6�&�
�"�h�G���P��� O��[��W���_�u�u�8��e����Où��Z�q\�� ��m�%�}�d�3�*����P���F��G1�*���f�m�%�u�j�)���&����P��F�X��1�"�!�u�~�W�W�������l ��W�����h�_�u�u�w�}��������EP��N�����!�%�f�
�"�n�E���Q���A��N�����u�u�u�u�'�2�(���J�ԓ�]ǻN�����d�3�
�a��l�K�������T��A�����0�<�0� �$�:��������l��h_�A���a�|�_�u�w�0�(�������9��R�����9�2�6�#�4�2�_�������U��Y�����4�
�:�&��+�C���?����u ��q(��Y���<�!�2�'�"�.����Q���F��G1�*���`�l�%�}�f�l��������O�d��Uʡ�%�c�
� �b�e����D�θ�C9��h��@���%�u�:�u�'�>��������  ��q(��3����|�_�u�w�0�(�������9��R�����9�
�
� �b�o����Hӂ��]��_����u�8�
�c�1��Oց�H���C9��[\��*���`�g�%�}�w�}�W������]ǻN�����b�3�
�d��n�K���&����lR��B1�L���}�d�1�"�#�}�F��Y����^��1��*��
�f�i�u�8�l����Aù��W��S�����d�n�u�u�#�-�@ށ�����l��S�����3�
�m�
�e�l�W������O��N�����3�
�a�
�e�a�WǪ�	����U��_��Fʴ�1�&�9�!�'����O����l�N�����3�
�f�
�f�a�W���&����P9��T��]���<�0� �&�0�8�_���&����e9��h]�*��y�g�|�_�w�}�;���K����_��X��*��� �d�d�
�d�a�W���Y�����V��M���-�3�
�m��n� ���Yە��l��\�� ��d�
�g�e�w�}�F�������9F�N��U���
�8�f�
�"�d�O���B�����O=�����
� �!�4�#�o�(���H����CT�
N�����2�6�#�6�8�u��������]9��E��*���x� �&�2�2�u�;���K����_��X��*��� �d�d�
�d�t�}���Y����A ��@1��*��
�f�i�u�w�}�W�������
9��hW�*��"�0�u�&�;�)��������9��^��H��r�u�9�0�]�}�W���Y����G��1��*��
�g�_�u�w�3��������G9��hW�*��i�u� �1�%�1� ���&����CU��X�����;�!�9�d�f�f��������l