-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ��m�d�a���(���
����GF�N�����9�u�u����;���:���F��h��U���������}���Y����G��T��;ʆ�����]�}�W�������	F��cN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�%�<���6����g"��x)��N���u�<�
�%�%�8���Cӯ��`2��{!��6�����u�f�w�2����I��ƹF��Y1�����
�u�u����;���:����g)��]����!�u�|�_�w�}��������G9��N��U���
���
��	�%���Hӂ��]��G�U���<�
�%�'�2�)�E��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����E�����u�u� �u���8���&����|4�_�����:�e�n�u�w�<�(�������\��b:��!�����
����_������\F��d��Uʴ�
�0� �;�e�g�8���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƭ�l��B��F��������4���:����U��S�����|�_�u�u�'�/����&����|3��d:��9�������w�n�W������]ǻN�����!�'�
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W�������\��yN��1�����|�_�9�f�}������P��RN�����:�u�g�m�f���������@FǻN�����4�!�4�
�8�.�(�������	F��s1��2���o�u�d�n�w�}��������R��X ��*���<�
�u�u���8���Y���A��N�����!�;�u�%���ށ�
����	F��s1��2������u�b�9� ���Y���F�^�D��u�u�6�;�#�3�W���*����9��Z1�Oʆ�������8���Lӂ��]��G��H���e�e�e�n�w�}��������R��c1��F���8�g�o����0���/����aF�
�����e�u�h�w�g�l�G��Y����\��V ������&�a�3�:�n�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���I����]ǻN�����4�!�4�
��.�B������5��h"��<������}�w�2����I����D��^�W�ߊu�u�:�&�6�)����-����l ��h[��U���
���
��	�%���Y����G	�N�U��e�e�w�_�w�}��������C9��Y����
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�e�w�]�}�W���
������T�����d�d�o����0���/����aF�
�����e�u�h�w�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�l�U�ԜY�Ư�]��Y�����;�!�9�d�g�g�$���5����l0��c!��]���:�;�:�e�w�`�U���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)����I����g"��x)��*�����}�u�8�3���Y���V�=N��U���&�4�!�4��2��������	F��s1��2������u�f�9� ���Y���F�L�U���6�;�!�;�w�-��������lW�=��*����
����u�W������F��L�W�ߊu�u�:�&�6�)��������_��h]��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��_�D��n�u�u�6�9�)����	����@��A]��F���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�D��e�w�_�u�w�2����Ӈ��P	��C1��F؊��o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��d�d�e�n�w�}��������R��X ��*���f�e�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�n�w�}��������R��X ��*���g�a�f�o���;���:����g)��_����!�u�|�o�w�m�G��H����D��N�����!�;�u�%�4�3����H¹�� F��d:��9�������w�l�W������F��L�E��d�e�d�n�w�}��������R��X ��*���g��o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�d�l�}�WϽ�����GF��h�����#�d�e�o���;���:����g)��_����!�u�|�o�w�m�G��I����]ǻN�����4�!�4�
�8�.�(���K����\��c*��:���
�����l��������\�_�D��d�d�e�n�w�}��������R��X ��*���g�f�u�u���8���&����|4�_�����:�e�u�h�u�m�G��H����]ǻN�����4�!�4�
�8�.�(���&����`2��{!��6�����u�`�3�*����P���V��^�N���u�6�;�!�9�}��������EP��N�&���������W������\F��T��W��d�e�n�u�w�>�����ƭ�l��D�����e�o�����4���:����S��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
����T��T��!�����
����_������\F��T��W��e�e�e�e�g�f�W�������R��V�����
�#�g�f�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����W��UךU���:�&�4�!�6�����&����F��d:��9�������w�k��������\�^�E��w�_�u�u�8�.��������]��[�*������o���;���:����g)��]����!�u�|�o�w�l�F��H����W��_�D��d�d�d�d�f�f�W�������R��V�����
�#�g���g�$���5����l0��c!��]��1�"�!�u�~�g�W��H����W��L�U���6�;�!�;�w�-��������9��q(��3�����u�u���8���&����|4�]�����:�e�u�h�u�l�F��H����W��_�D��d�d�d�d�f�l�F��H����W��_�D��u�u�6�;�#�3�W�������l
��1��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�D��w�_�u�u�8�.��������]��[�*��o������!���6���F��@ ��U���o�u�e�e�g�l�G��[���F��Y�����%�6�;�!�;�l�(��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��_�E��n�_�u�u�>�3�Ͽ�&����@�=��*����
����u�W������F��L�E��w�_�u�u�#�/����Y����V��S��U���!�<�2�_�w�}��������U��R �����u�3�4�
��;���
����_F��L�����_�u�u�<�9�1��������V��c1��D���8�e�o����0���s���@��V�����2�7�1�g�w�}�8���8��ƹF��^	��ʴ�
�<�
�&�&��(���&����F��d:��9����_�u�u�>�3�Ͽ�&����Q��V��U�����n�u�w�.����Y����U��\��D��������4���Y����W	��C��\�ߊu�u�<�;�;�;�(�������^9��h��*��a�o�����4���:����U��S�����|�_�u�u�>�3�Ϸ�&����\��X��Dۊ� �g�e�%�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������9��h(��*���%�d�
�0��l�E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V�����&�$��
�#�����Y�Ɵ�w9��p'�����u�<�;�9�6���������\��x!��4��u�u�&�2�6�}��������lT��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2���������Q�=��*����
����u�W������]ǻN�����9�0�<�6�9����M����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�g�1��Bׁ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�
�0��l�B��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��Q=��8���,� �
�f�1��Fׁ�K����g"��x)��*�����}�d�3�*����P���F��P ��U���-� ���#�o�(���&����\��c*��:���
�����l��������l�N�����u�&�0�
�2��F��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*���
�&�$���)�(���&����`2��{!��6�ߊu�u�<�;�;�<�(���&����
R�,��9���n�u�u�&�0�<�W���&�Փ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������_��N��1��������}�B�������V�=N��U���;�9�!�%�f����K����	F��s1��2������u�g�9� ���Y����F�D�����8�
�l�'�0�l�N���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��(�����a�
�g�o���;���:����g)��_����!�u�|�_�w�}����Ӡ��A��\�U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_�������V�=N��U���;�9�!�%�e�����K���5��h"��<������}�w�2����I��ƹF��^	��ʼ�8�b�3�
�`��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��^��B���2�d�d�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lP��Q��LҊ�f�o�����4���:����S��X����n�u�u�&�0�<�W���&�֓�V��\�Oʆ�������8���Lӂ��]��G�U���&�2�4�u��<�E�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�
�6�o�B�������
F��d:��9�������w�n�W������]ǻN�����9�4�
�<��.����&����U��N�&������_�w�}����Ӈ��@��U
��D��o�����W�W���������D�����'�2�d�f�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������l��h_�E��������4���Y����\��XN�N���u�&�2�4�w�8����&����@9��hW�*��o������!���6�����Y��E��u�u�&�2�6�}��������A	��E��D��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1�%���¹��_9��R��*���b�3�
�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��Y	��*���
�;�&�g�>�l�(���&����\��c*��:���
�����}�������9F������4�'�9�
�8�����Hʹ��V9��1��*��c�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Z��D��&���!�
�&�
�w�}�#���6����9F������4�
�<�
�3��D���Y����v'��=N��U���;�9�4�'�;���������
9��R1��F���
�e�e�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����R��[�����:�%�d�
���(ځ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�'��)�1���5����_��h��*ۊ� �d�m�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��3����:�
�l�e�8�F�������
^��N�&���������W��Y����G	�UךU���<�;�9�4�%�1�(���&����lW��1��D���3�
�d�g�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h'��0����0�8�a���(���&����	F��s1��2������u�d�}�������9F������6�
��������Mǹ��9��P1�C��������4���Y����W	��C��\�ߊu�u�<�;�;�<����&����	��h_��G���e�c�'�2�f�e�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�����'��:�
�n�o��������V�=��*����
����u�FϺ�����O��N�����4�u�9����%�������l��h��*��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���0����r4��R��A܊�
�
�0�
�n�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��3����:�
�
�2��G���Y����)��t1��6���u�d�1�"�#�}�^�ԜY�ƿ�T���������!�g��(�E���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�
���,�"��D���&����CW�=��*����
����u�FϺ�����O��N�����4�u�'�
�"�o�E���Y�Ɵ�w9��p'��#����u�c�u�8�3���B�����Y�����&�2�
� �e�h����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����%�
� �g�e�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��S1�����
� �g�`�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��R	��*���f�m�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ʃ�C9��G1�����g�
�a�o���;���:����g)��_����!�u�|�_�w�}����Ӓ��lR��Q��D؊�d�o�����4���:����P��S�����|�_�u�u�>�3�Ϫ�	����F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��n����NŹ��\��c*��:���
�����l��������l�N�����u�8�
�l�1��Oׁ�H����g"��x)��*�����}�u�8�3���B�����Y�����f�
� �f�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h�����l�
�g�o���;���:����g)��[�����:�e�n�u�w�.����Y����^��B1�C���u�u��
���(���-���T��X����n�u�u�&�0�<�W�������lW��Q��Dي�d�o�����4���:����S��S�����|�_�u�u�>�3�ϳ�����l ��_�����u��
����2���+������Y��E��u�u�&�2�6�}����I����U��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�o�(���M�ӓ�F��d:��9�������w�l�W������]ǻN�����9��
�
�"�i�G���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y������3�
�g��n�Mύ�=����z%��r-��'���f�1�"�!�w�t�}���Y����R
��Z��@���
�c�
�a�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��h��A���%�u�u����>���<����N��
�����e�n�u�u�$�:����K�ԓ�R��Q��A݊�d�o�����4���:����U��S�����|�_�u�u�>�3�Ϸ�����lR��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��A���&����CT�=��*����
����u�FϺ�����O��N�����4�u�8�
�`�;�(��&���5��h"��<������}�d�9� ���Y����F�D�����8�
�m�3��d�(��Cӵ��l*��~-��0����}�f�1� �)�W���s���@��V�����a�3�
�`��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���`�d�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƿ�\��R��*���`�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��@���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l��C1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������9��h[�*��o������!���6�����Y��E��u�u�&�2�6�}����N����U��G]��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�k�(���L�ߓ�F��d:��9�������w�h�W������]ǻN�����9�!�%�c��(�B���	����`2��{!��6�����u�`�w�2����I��ƹF��^	��ʡ�%�c�
� �b�e����Y����)��t1��6���u�`�u�:�9�2�G��Y����Z��[N��'���9�
�
� �b�i����Y����)��t1��6���u�`�u�:�9�2�G��Y����Z��[N����
� �`�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������V��F���
�d�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������^��1��*��
�d�o����0���/����aF�
�����e�n�u�u�$�:����&����P��N�&���������W������\F��d��Uʦ�2�4�u�
�����J����	F��s1��2������u�g�9� ���Y����F�D�����7�3�
�a��n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h�����d�3�
�l��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���c�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�e��hZ�� ��l�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Q��B1�@���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Oƹ��lS��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2���������9��T��!�����
����_�������V�=N��U���;�9�!�%�1��Cށ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�e�3��i�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�
� �c�n�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��D�����a�1�8�'�6����H����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�d��(�A���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʦ�:�0�0�2�����J����	F��s1��2������u�d�}�������9F������!�%�f�
�"�k�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����3�
�m�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������
9��hY�*��o������!���6�����Y��E��u�u�&�2�6�}��������U��[��D��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����P��N�&���������W��Y����G	�UךU���<�;�9�!�'�i�(���N�֓�F��d:��9�������w�h�W������]ǻN�����9�9�
� �`�k����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���b�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ�� T��B1�E���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����N¹��lQ��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��C���&����CT�=��*����
����u�W������]ǻN�����9�'�#�
�"�j�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����6�&�
� �a�i����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N����
� �b�m�'�}�W���&����p9��t:��U���u�:�;�:�g�f�W���
����_F��Y	��*���
� �b�g�'�}�W���&����p9��t:��U���u�:�;�:�g�f�W���
����_F��a1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������]��h�� ��g�%�u�u���8���&����|4�N�����u�|�_�u�w�4����+����9��[1����� �b�a�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������R��1�����0�
�
�
�"�e�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����d�4�9�:�2��(���N�Г�F��d:��9�������w�m��������l�N�����u�8�
�c�1��E߁�K����g"��x)��*�����}�u�8�3���B�����Y��'���0�
�9�
�2�2�(���A�Г�F��d:��9�������w�m��������l�N�����u�4�2�d�6�1����
�ד�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Cہ�����l^��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��O���&����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�n����O����\��c*��:���
�����}�������9F������&�9�!�%�c�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʺ�
�:�1�f�>�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʇ�;�0�
�9��3����&����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�h����Nǹ��\��c*��:���
�����}�������9F������%�l�
�
�"�e�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V��*���<�3�
�f��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�l�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����P��N1�����
�b�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�g�<�3��e�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
�9�
�0�8��(�������l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�o�(���@�ӓ�F��d:��9�������w�m��������l�N�����u�8�f�
�"�d�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�g�
� �n�m����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���3�
�g�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��M���
�f�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�CU��Q��@؊�g�o�����4���:����V��X����n�u�u�&�0�<�W�������D9��hW�*��o������!���6�����Y��E��u�u�&�2�6�}�(�������T��^1��*���
�g�o����0���/����aF�
�����e�n�u�u�$�:��������_	��Y�����c�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����l��X�����;�!�3�
�`��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��U�����<�<�;�!�1��Aׁ�K����g"��x)��*�����}�u�8�3���B�����Y�����`�
� �l�d�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E����� �l�e�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���d�e�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G]�����e�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӗ��R
��1�����
�m�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������V
��Z�*���l�m�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƹ�l��x��Fӊ�:�4�
�
�"�l�Fف�J����g"��x)��*�����}�d�3�*����P���F��P ��U���-� �,� ��(��������U��\�����u��
����2���+������Y��E��u�u�&�2�6�}��������l*��G1�*ڊ�
�
� �d�e��C��*����|!��h8��!���}�e�1�"�#�}�^�ԜY�ƿ�T����*����'��:��d�G���I�ԓ�F9��W��D��������4���Y����W	��C��\�ߊu�u�<�;�;�<����&����	��h_��G���e�3�
�e�n�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�f��(���&����lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���?����\	��W��*���
� �d�a��o�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�����'��:�
�n�o����K����V��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�6�/��������\��1�����a�3�
�d�b�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����g�
�0�o���;���:���F��P ��U���'�!�'�
��/���*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��^	��ʴ�
�0� �;�f�-����Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�D�����%�'�!�'������Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������4�
�0� �9�n����Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����u�%�'�!�%��(�������g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����9�4�
�0�"�3�B�������`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����4�u�%���.�W���-����t/��a+��:���`�1�"�!�w�t�}���YӅ��C	��Y��G��d��3�e�1�(�(���
����@9��h_�����&�u��u�w�:������ƹF�N��1������]�}�W���Y����`2��rN�<�����_�u�w�}�W���I����g.�'��0���n�u�u�u�w�9�ށ�0����	F��c+��'�ߊu�u�u�u�8�)� ���1����}2��r<��N���u�%�'�u�]�}�W���Y����\��yN��1��������}�D�������V�=N��U���u�<�d�o��}�#���6����e#��x<��F���:�;�:�e�l�}�W���Yӂ��GF��x;��&���������W��Y����G	�N����u�;�u�:�'�3���s�����G�����g�m�d��1�m��������]��1�<�ߊu�u�0�0�>�}�}���Y���z"�'��0���n�u�u�u�w��:���8���/��r)��N���u�u�u�1�9��>���Y�ƅ�g#��eUךU���u�u�:�!� ��?��0����v4�d��Uʥ�'�u�_�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u�%�.���0�Ɵ�w9��p'�����u�u�u�<�g�g�>���-����t/��a+��:���c�u�:�;�8�m�L���Y�����N��U���
���n�w�}�W�������	F��cN��1��������}�D�������V�UךU���;�u�:�%�9�3�L�ԶY����\��Y��U���m�d��3�g�;����J����R��'��U���2�;�'�6��}�W���Yӯ��	F��c+��'�ߊu�u�u�u���#���Y�ƅ�g#��eUךU���u�u�<�e� ��?��0����v4��N��U���1� �
���}�W���<����]ǻN�����}�u�u�u�w�9����Y����g"��x)��*�����}�d�3�*����P���F�N�� ���u� �u����>���<����N��
�����e�u�n�u�w�8�Ͻ�����]��=d�����_�u�u�
��0�������]��1�����1�%� �u�w�2�����ơ�w^��*��*ڊ�8�9�f�;��o���&¹��K9��Gd��Uʲ�;�'�6�8�'�u�W���Y����wF�_�U���u�u�����2��Y��ƹF�N��������h�w�o�}���Y���W��h9��!���k�f�y�u�w�}�WϺ�����w2��
P��G�ߊu�u�:�!�:�-�_���Y�����N��U���-� ���#�o�(���K�ޓ�JǻN��U���<�d�h�u��%�"���6���� 9��h\�*��_�u�u�u�w�2���Y����~3��N!��*���3�
�d�
�e�f�}���Y����@��Q��A���f�
�
�d�w�}��������^T��_��A���
�<�:�%�a�3�(���K�����R��U���u�_�u�u�w�}�3��Y��ƹF�N�� �����u�k�e�W�W���Y�ƨ�]V��~*��U��c�y�u�u�w�}����&����{F�]����u�:�!�8�'�u�W���Y����_�	N��*���y�u�u�u�w�/����D�ƭ�l��d��U���u�1�;�u�i�:����&����CV�N��U���6�u�k�2�'�;�(��&����F�N�����u�k�2�%�1��E݁�H��ƓF�Q1�����!�f�;�
�c�l�"��CӅ��C	��Y��G��d��3�e�1�8�������lWǻN�����<�u�4�u�]�}�W���Y���F��=N��U���u� �
���}�I��s���F�S��*����u�k�f�{�}�W���Yӂ��G9��s:��H���a�_�u�u�8�)����Q���F�
��E��u�
�&�<�9�;�(��&����F�N�����u�k�1�4�$�:�(���K�ӓ�O��=dװ���u�x�!�0�4�/����
����N��h-�����u�3�!�0�$�<�ϳ�����F�=N��U����
�&�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���	����U��S�����
�!�
�&��f�W���Y���F��[��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����s���F�N��U���u�u�4�
��;���Y����`9��ZUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W������G��h^�����4�&�2�u�%�>���T���F��h�� ���e�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���	����F��1�����h�4�
�:�$�����I���F�N��Uʰ�&�_�u�u�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C]�����|�4�1�;�#�u��������F9��1��U���%�6�;�!�;�l�G���PӒ��]FǻN��U���u�u�u�u�w�}��������9��R	��Hʴ�'�9�
�:��2���&����9��E��D��_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����E�����
�'�2�4�$�:�W�������K��N�����0� �;�d�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���R��R�����%�0�u�h�6�����&����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9����Q����P	��h��G���%�u�u�%�4�3����H���O��_�����u�u�u�u�w�}�W���Y����V��Y1�����u�h�4�'�;���������
9��R1�����d�e�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F������'�
�
�'�0�<����Y����V��C�U���4�
�0� �9�o����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�V�����;�g�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�������V��T��*���g�a�%�u�w�-��������lV�G�����_�u�u�u�w�}�W���Y���R��R�����%�0�u�h�4��9���8����A��1��E���2�d�c�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C�����!�'�
�
�%�:�����Ƽ�\��D@��X���u�4�
�0�"�3�D�������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��*��� �;�f�%�2�}�JϿ�&����G9��\��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ�ӈ��N��^����� �g�a�%�w�}��������EW��G��U���;�_�u�u�w�}�W���Y���F��h�� ���f�%�0�u�j�>�(���<����G��hZ�����'�2�d�g�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���'�!�'�
��/�Ͽ�
����C��R��U���u�u�4�
�2�(����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N�����0� �;�a�'�8�W������]��[�*��u�u�u�u�w�}����s���F�N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!��.�(�������\�R�����
� �g�a�'�}�W�������l
��h^��\���=�;�_�u�w�}�W���Y���F�V�����;�a�%�0�w�`����7����a4��E��C���e�'�2�d�c�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���%�'�!�'����������]F��X�����x�u�u�4��8����L����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʴ�
�0� �;�b�-����DӇ��P	��C1��F؊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�����PӇ����F�����;�
� �g�c�-�W���	����@��A_��\���u�=�;�_�w�}�W���Y���F�N��*��� �;�`�%�2�}�JϽ�&����k'��C��*���0�d�'�2�f�i�}���Y���F�N�����<�n�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=d��U���u��9�
�8�����
����lT�������%�:�0�&�w�p�W�������l ��h"�����'�2�g�c�6�.���������T��U´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������W������u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���u�u�u�u�>���������C9��E��G��i�u��9��2�(���	����A��_�N���u�u�u�u�w�}�Wϻ�
�����T�����2�6�d�h�6�����
����g9��1����|�!�0�u�w�}�W���Y���F�N��9���
�:�
�:�'�.����K���F��h�����#�
�n�u�w�}�W���Y����������u�u�u�u�w�3�W���Y���F���U���_�u�u�;�w�/����B���F������%�:�0�&�w�p�W���	����@�V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���H����[��N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�(���&�����Yd��U���u�u�u�u�w��(���&����Z�q\�� ��m�%�n�u�w�}�W���Y�����GY�����g�l�i�u�4�-�(���J�֓�]ǻN��U���u�u�u�u�$�8�(���&����Z�^��*��� �f�m�%��n��������]ǻN��U���u�u�u�u�:��N�������F���*���3�
�a�
�e�W�W���Y���F�N����
�0�
�g�e�a�W���&�ԓ�F9��1��N���u�u�u�u�w�}�WϪ�	����A��_�U��!�%�`�
�"�n�O���B���F�N��U���u�8�
�e�%�:�F��Y����^��1��*��
�f�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=N��U���4�&�2�u�%�>���T���F��X�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������A��N���ߊu�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�ӓ�@��G�����_�u�u�u�w�}�W���Y����VW��[�����g�<�d�
�2��E��E�ƞ�]��h��*���&�g�<�d��(�N���	��ƹF�N��U���u�u�0�0�2�����&����T��R�����!�1�/�'�$�;�(��&����F�N��U���u�u�;�"�>�3�������� S�
N��#���
�
� �c�a�-�_������\F��UךU���u�u�u�u�w�}�(���K�ӓ�V��\�I���
�4�g�`�1��Aف�J���F�N��U���u�!�%�f��8�(��I���G��W�� ��c�%�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�&�<�;�'�2����Y��ƹF��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G��U���;�u�u�u�w�}�W���YӇ��l
��q��9���
�l�g�0�g�k����H���F��E1��*���
�:�%�d���(߁�&����Q��G]�U���u�u�u�u�w�}��������A9��X��L���0�d�'�2�f�m�K�������l ��h"����
�
�
�
��(�F��&����F�N��U���u�u�6�
���6�������9��1����c�i�u�'��)�1���5����_��h��*ي� �d�b�
�d�W�W���Y���F�N��*������0�:�i�(���&����^��S�����!��'��8��N����ד�l ��^�*��_�u�u�u�w�}�W���Y����}"��v<�����a�
�
�
�2��D���DӇ��l
��q��9���
�l�g�0�g�l����I�Г� ]ǻN��U���u�u�u�u�;��3���+����^9��h��*���
�l�u�h�6�/��������\��1�����`�3�
�d�e�-�L���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�u�u�x�w�.����	����@�CךU���'�6�&�u�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H��r�u�=�;�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�����d�|�u�=�9�}�W���Y���F������
�0�8�l��8�(��M���T��Q��G؊�d�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǻN��Xʴ�&�2�u�'�4�.�Y��s���C��R��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������A�C�����u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���J����lT�V ��]���!�:�1�3��n�(��DӇ��P	��C1��D��|�u�=�;�w�}�W���Y���F��d1�� ����!�g�
�2��F��E�ƪ�l��{:�� ���f�3�
�d��o�}���Y���F�N�����!�%�
�0��l�B��Y����G��h��G���%�n�u�u�w�}�W���Y����V
��Z�����d�b�i�u�2���������l��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}���Y���R��P �����&�{�x�_�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�f�1�0�E���Y����9F�N��U���u�u�u��;���������9��P1�@���h�<�
�<��/�;���&�ד�F9��1��N���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B���F���U���!�&�4�0��-�9���
����UF��RN�����8�6�<�0�w�p�W�������l ��h�����%�:�u�u�%�>��������R����6���&�y�4�
�2�}��������F9��1��\���u�7�2�;�w�}�W�������R��d1��ʼ�_�u�u�u�w�}�W���Ӈ��`2��C_�����u�k�_�u�w�}�W���Y���Z �F��*���&�
�:�<��}�W�������]��X�����!�'�u�u�'�>��������lV�G�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�e�;���s���F�N��U���0�&�_�u�w�}�W���Y���F�V��&���8�i�u�%���ށ�
����9F�N��U���u�u�u�;�w�;�}���Y���F�@��U����
�!�
�$��W���s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�D�������F�N��U���u�u�0�&�]�}�W���Y���F�N������3�8�i�w�-�$�������^9��=N��U���u�u�u�u�w�3�W���s���F�N�����u�%��
�#�����Y���F�N��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�8�u��������U��Z��G��4�
�:�&��+�(���P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y���F��[��U���4�
�:�&��2����Y�ƭ�l����U°�<�6�;�
�"�o�C���Y�ƭ�l��D��ۊ�|�|�!�0�]�}�W���Y���F�N������3�8�i�w�-�$���ǹ��^9��=N��U���u�u�u�u�w�1����Y���F�N��U���u�%��
�$�}�JϿ�&����GU��D��N���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�=�;�4��	��������[�=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���4�
��3�:�a�W���*����9��Z1����u�u�u�u�w�}�W������F�N��U���u�u�u�%������DӇ��`2��CZ�����n�u�u�u�w�}�W���YӃ����=N��U���u�u�u�=�9�<�(���
�ӓ�@��S����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�4�
��;���Y����g9��1�����_�u�u�u�w�}�W���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:��ߊ�&�
�n�u�w�}�W���Y����������u�u�u�u�w�5�Ͽ�&����GP��D��U��_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�6��$������R��c1��F���8�g�_�u�w�}�W���Y���V
��=N��U���u�u�u�u�w�}�W���7����^F���&���!�
�&�
�l�}�W���Y���F���U���_�u�u�u�w�}�W���Ӊ��V��
P�����u�u�u�u�w�}�W���7����^F�L��-���w�_�u�u�w�}��������F�R �����0�&�_�u�w�}�W���K����G9��hZ�*��i�u�!�
�8�4�(�������V��RF�����}�g�g�3��i�(��U���lǻN��G���3�
�a�
�d�a�W���Y��� ��E��D��u�=�;�}�:��G���&����CT�N��R��u�9�0�_�w�}�W�������l ��]����u�u��
�"�n�O���Y����G��X	��*���!�'� �&�0�8�_�������l
��1�F���u�;�<�;�3�)��������9��G�U����;�0�
�;�����H����R��G\��H���8�f�
� �`�m�����Ƹ�C9��h��B���%�|�_�u�w�<��������]��1��D݊� �l�a�%�w�`�_�������Z9��hX�*��4�1��;�2���������l��B1�G���|�_�u�u�6�:�F�������@9��^1��*��
�f�i�u�w�}�W���+����9��[1����� �m�a�%�w�5��������W_��^1��*��
�g�e�u�w�l�^ϻ�
��ƹF�N�����8�g�
� �o�i���Y����R��1�����0�
� �m�c�-�W��Q����VT��[�����d�<�3�
�g��DϿ�Ӵ��T��V�����
�
� �b�a�-�^�ԜY�ƞ�]��h��*���:�
�
� �o�i����D������YN�����
� �a�f�'�}�W�������l
��1�U���0�w�w�_�w�}����H����l��X��*��� �m�m�%�w�`�}���Y���C9��h�� ��g�%�u�=�9�u��������Z9��hV�*��e�u�u�d�~�8����Y���F��R����
� �m�e�'�f�W���+����9��[1�����3�
�g�
�e�a�Wǌ�����R
��X ��*ۊ� �b�c�%�w�2�W�������l
��h_����u�4�2�g��l����A����Z�D�����6�#�6�:��5��������F��P ��]���
�
� �a�d�-�^ê�&����T��B �����}�e�u�u�:��B���&����CW�C����!�u�|�|�~�W�W�������l��h�����<�3�
�e��n�K���Y���F��V ��G���9�:�0�
�"�j�C���Y����N��h�����<�3�
�b��o�G���Y�����RNךU���u�u�0�d�1��A߁�K���F��Y	��*���
�;�&�3��d�(��E���F��R ��'���0�
�
�
�"�j�E���Y�ƾ�e9��hY�*��u�9�0�w�u�W�W���T�ƭ�l��RN�����u�'�6�&�y�p�}���Y����\��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����VJ��G1�����0�
��&�d�;���Y����P	��h��G���%�|�u�u�5�:����Y�����F�����4�
�:�&��2����Y�ƭ�l��E��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^�������C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*���� 9��Z1�U���u�:�}�0�>�>��������l��
N��*���&�
�#�
�~�t�^Ϫ���ƹF�N��U���%�1�;�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��X ��I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���0�4�&�2�w�/����W���F�V�����4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�N�����;�u�u�u�w�4�W�������C9��Y�����6�d�h�4��)����Y������T�����2�6�d�h�6�����
����g9��1����|�u�=�;�]�}�W���Y���R��S��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�<�(������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������R��V�����'�6�&�{�z�W�W���	����W��D�����:�u�u�'�4�.�_�������C9��P1������&�f�3�:�o�W�������l ��]�����u�u�7�2�9�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1����u�;�u�:��8��������lT��h�Hʴ�
�:�&�
�!��^���Y����l�N��U���u�4�
�0�3�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���%�'�!�'��}����Ӗ��P��N����u�%�'�!�%��(�������A	��N�����&�4�
�0�w�-��������`2��C]�����y�0�<�6�9����M������h��3����:�
�l�e�8�G�������^�V�����;�e�%�0�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�f�3�8�e�}��������K��X �����f�
�g�h�6�����&����O�N�����u�u�u�u�w�}��������lV�
N�����
�:�
�:�'�l�(݁�&ù��A��[����u�u�u�9�2�W�W���Y���F��h�� ���e�i�u�%�%�)����&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�0� �9�l�����Ƽ�\��D@��X���u�4�
�0�"�3�F���
����C��T�����&�}�%�6�{�<�(���&����l5��D�����g�u�-�!�8�9����Jǹ��F��E1��*���
�:�%�d���(ށ�����J��G1�����
�
�'�2�]�}�W������F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<�ϰ��Ω�Z��Y
�� ��a�%�u�u�'�>�����ד�O����ߊu�u�u�u�w�}��������F���*����'��:��d�E���H����lW��d��U���u�0�&�u�w�}�W���Y����C9��C��*���h�4�
�0�"�3�F�����ƹF�N�����3�u�u�u�2�9��������9l�N�U���'�!�'�
�w�.����	����@�CךU���%�'�!�'����������PF��G�����4�
�0�u�'�.��������l��h��*���0�<�6�;��(�E���	����_9��s+��'���'�
�a�0�g�/���O�ƭ�l��B��G���0�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��F���8�g�u�;�w�2�_ǻ�����W9��h\�*��h�4�
�:�$��ށ�P���G��d��U���u�u�u�4��8����K���P
��y*��4���0�8�a�
������M��ƹF�N�����_�u�u�u�w�}�W�������]9��S�����!�'�
�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h�� ���f�4�&�2�w�/����W���F�V�����;�f�4�&�0�����CӖ��P�������4�
�<�
�$�,�$�������^9�������1�3�
�f��o�W���0����r4��R��Aފ�
�
�0�
�o�q��������lU��E�����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GU��D��\ʴ�1�;�!�}�/�)��������9��S�����;�!�9�d�g�t�^Ϫ���ƹF�N��U���%�'�!�'��}�JϽ�&����k'��C��*���0�d�'�2�f�o�}���Y���V
��d��U���u�u�u�4��8����J���R��R�����%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������G��hZ�����;�%�:�0�$�}�Z���YӇ��A��E ��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�n����K�Ʃ�Z��Y
�� ��a�%�y�6���2���+����lR��R1�����d�a�u�%�%�)����&����l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����0�<�6�;��(�E���	���R��X ��*���
�|�|�u�?�3�}���Y���F�V�����;�a�i�u�;��3���+����^9��h��*���
�f�n�u�w�}�Wϻ�
��ƹF�N��U���%�'�!�'��}�JϿ�&����A��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������R��P �����&�{�x�_�w�}��������9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�
�&��q��������U��Z��G���9�����)����O����l��h_�Yʴ�
�0� �;�b�-����Y����V��=N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�d�;���Y����]	�������1�3�
�f��o�JϿ�&����G9��1�\���!�0�u�u�w�}�W���YӇ��A��E ��U��6�
��������MŹ��9��P1�A�ߊu�u�u�u�;�8�}���Y���F�V�����;�`�i�u�'�/����&ƹ��V��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h_�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�a�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h_�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�`�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(������]F��X�����x�u�u�4��4�(���&�ғ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��N�U´�
��3�8�g�9� ���Y�����T�����d�d�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�h�W�������A	��D�X�ߊu�u�%�&�0�?���&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����^�
N�����;�!�9�d�f�`����*����W��X����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�c�<����Y����V��C�U���4�
�<�
�3��C���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������[�V�����
�#�
�u�w�-�4���
����W	��C��\��u�u�0�1�'�2����s���F������7�1�l�u�$�4�Ϯ�����F�=N��U���&�2�7�1�n���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����M�����T�����d�d�h�4������Jӂ��]��G����u�;�u�'�4�.�L�ԶY���F��h��*���$��
�!��.�(���
������T��[���_�u�u�%�$�:����&����GW��D��*���<�;�%�:�w�}����
�έ�l��h��*��_�u�u�0�>�W�W���Y�ƥ�N��h��*���
�a�u�=�9�W�W���Y���F��h��*���$��
�!��.�(���DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����<�
�&�$���ށ�
����[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�ƭ�l��h�����
�!�
�&��}����Ӗ��P��N����u�%�&�2�4�8�(���
�ԓ�@��h�����%�:�u�u�%�>����	����l��h[����u�0�<�_�w�}�W����έ�l��h��*��u�=�;�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��F1��*���
�&�
�u�$�4�Ϯ�����F�=N��U���&�2�6�0��	��������l��^	�����u�u�'�6�$�u��������lQ��=N��U���<�_�u�u�w�}����	����l��hY�U���;�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������B9��h��*���
�u�&�<�9�-����
���9F������6�0�
��$�i����J����Z��G��U���'�6�&�}�'�.��������9F����ߊu�u�u�u�1�u��������l_�����ߊu�u�u�u�w�}��������B9��h��*���
�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����Z��D��&���!�
�&�
�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�.��������l��h��*���&�<�;�%�8�8����T�����D�����
��&�`�1�0�C���
����C��T�����&�}�%�&�0�?���O���F��P��U���u�u�<�u�6���������O��_�����u�u�u�u�w�-��������`2��C[�����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GP��D��U���<�;�%�:�2�.�W��Y����C9��P1������&�c�3�:�h��������\������}�%�&�2�5�9�F��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��h��*���h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���
����@��d:��܊�&�
�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���'�
�!��%�����@�֓�lV��h��D��
�d�i�u�#�����&����\��R�� �&�2�0�}�%���������C9��h^��*ڊ� �d�g�
�c�q�E���s���R��[�����:�%�d�
���(���H����CR�
N��*�����!��5�/����O����V��h�F���:�;�:�d�l�}�WϿ�����u	��{��*���e�0�d�3��m�D���Y����G��X	��*���!�'� �&�0�8�_���&����\��X��Dӊ�
�
�
�
�"�l�Dց�H���F��P ��]���-� �,� ��(��������U��\�����n�u�u�4�%�1�(���&����lW��1��E���3�
�e�c�'�}�J�ԜY���F��h'��0����0�8�a���(���&����D��F�����%�
�0�
�f�h�G���Y�����RNךU���u�u�'�
�#���������lT��h^�� ��a�
�f�_�w�}��������l*��G1�*؊�
�
�
� �f�k�(��E��ƹF�N�����!��'��8��N����֓�l ��^�*��"�0�u�&�;�)��������N��S��D���0�&�u�u�w�}�WϽ�&����k'��C��*���0�e�'�2�f�k�}���Y����_��X�����d�
�
�
�����Nù��Z�=N��U���u�9��������&�ғ�lV��R	��A���=�;�}�0��0�E�������N��S��D���0�&�u�u�w�}�WϿ�����u	��{��*���g�0�e�g�1��G���	��ƹF��E�����'��:�
�n�o����L����V��h�I���u�u�u�u�6�/��������\��1�����g�3�
�e�n�-�W����ο�_9��G\�����d�`�e�u�w�l�^ϻ�
��ƹF�N�����!��'��8��N����֓�l��h_�N���u�4�'�9��2�(���	����9��1��*��l�%�u�h�]�}�W���Y����}"��v<�����a�
�
�
�2��D������@��C�����d�`�}�|�j�z�P������F�N�����9�
�:�
�8�-�Fց�&����9��h_�L���n�u�u�4�%�1�(���&����lW��1��D���3�
�e�a�'�}�J�ԜY���F��E1��*���
�:�%�d���(ށ����� 9�������0�
�8�g�%�:�F��Q���A��N�����u�u�u�u�6�/��������\��1�����'�2�d�e�]�}�W���&����\��X��Dӊ�
�
�
�
�"�l�Nށ�J���9F�N��U���
�!��'��2�(���I����l ��^�*��"�0�u�&�;�)��������N��S��D���0�&�u�u�w�}�WϽ�&����k'��C��*���0�d�'�2�f�o�}���Y����_��X�����d�
�
�
�����@˹��Z�=N��U���u�9��������&�ғ�lW��R	��M���=�;�}�0��0�E�������N��S��D���0�&�u�u�w�}�WϿ�����u	��{��*���g�0�d�g�1��G���	��ƹF��E�����'��:�
�n�o����M����W��h�I���u�u�u�u�4��9���8����A��1��D���2�d�a�"�2�}��������V��[�E���u�d�|�0�$�}�W���Y����A��C1�����:�
�l�e�2�l����I�Փ�]ǻN�����!��'��8��N����ד�l ��_�*��i�u�u�u�w�}����7����a4��E��C���d�'�2�d�c�*����
����^��E��D��}�|�h�r�p�}����s���F�V�����:�
�:�%�f��(���&ǹ��lW��1��N���u�7�8�'�2�;�(��&���F��Y
�����
�:�
� �n�o����Ӗ��9��Z�����
�:�
� �n�i����s���Q��E	�����;�!�3�
�a��E��Yۖ��9��Z�����
� �l�b�'�}��������_	��Y�����c�
�g�n�w�}���� �ד�l ��Y�����h�}�0�
�:�l�(���O�ѓ�F��SN����
� �c�f�'�t�}���Y����@��h��G���%�u�h�3���;�������l��h_�@�ߊu�u�0�0�2�����&����P��N�U���u�u�u��9�8�(���&����lT��h��M���%�u�=�;��<����&����lP��h�E���u�d�|�0�$�}�W���Y����R��1�����'�&�g�<�1��Nׁ�J���F��^����� �g�a�%�w�`�U���������[�����:�%�&�'�0�o�A������]��[��F���9�0�w�w�]�}�W���&����e9��h]�*��i�u�'�2��;�(��&���F��@ ��U��n�u�u�3���;�������l ��_�����h�3�
�:�2�)����I����lW��UךU����-� ���)�E܁�����l��S��U���u�u�<�
�'�/����Iӑ��]F��R�����3�
�`�
�e�m�W���H����_��=N��U���u�0�
�8�f�;�(��&����9F�C����3�
�g�
�2�<����Y����V��C�U���2�%�3�
�e�����
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�y�4��8�W���
����@��d:��؊�&�
�|�u�w�?����Y���F��QN��]���6�;�!�9�0�>�F������F��SN��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�W���Qۇ��@��CN�����:�&�
�:�>��^�������C9��Y�����6�d�h�4��4�(�������@��Q��D���|�!�0�u�w�}�W���Y����A��B1�G���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W�������lT��h��I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B���F��G1��*��
�e�i�u�#�����&����\��R�� �&�2�0�}�9�����&���O�=N��U���9�
�:�
�8�-�Fށ�����l��S�����:�<�
�0�#�/��������Z*��^1�����:�
�
�0��m�^�������]��V�����
�#�
�|�l�}�WϷ��ѓ�F9��1��U��w�w�"�0�w�.����Q����^��B1�E���|�k�&�2�2�u��������EW��G�����u�e�n�u�w�4��������l��S��D���=�;�}�8��h����O¹��[��G1�����9�b�e�u�;�8�U���s���Z��h8�� ��m�%�u�h�3�<����&����S��UךU����3�
�f��l�K�������l �� ]�����u�u�u�:�9�2�G��Y����R��h_�� ��b�%�u�h�$�9��������G	��B �����}�%�6�;�#�1�Bہ�P����]��Y�����&�9�
�f�1��F܁�H����F�Z��#���
�g�
�f�k�}�W���Y����R��h_�� ��b�%�u�=�9�u����&����W��^��H��r�u�9�0�]�}�W���Y����@��h_�����d�
�d�_�w�}��������Z9��hY�*��i�u�!�%�c����O����R��E��*���b�e�%�|�]�}�W������� 9��Q��EҊ�g�i�u�!�'�i�(���N�Г�F��SN�����
�g�
�g�l�}�WϮ�@ƹ��U��^��G��u��;�0��1�(�������U��Z��Gʺ�u�0�
� �`�m����s���C9��h
�����;�<�3�
�b��E��Yے�� R��B1�G���u�'�1�9�#�9����
����lW��G�U���%�l�
�0�8�:��������F9��1��U��}�
�b�1�:�/����&����Q��N��ʴ�
�:�&�
�!��^�ԜY�Ƽ�
^��h��M���%�u�h�}�:��A���&����CT��Y
�����d�4�9�/�%�.����KŹ��]ǻN��*��� �!�d�
�"�i�D���Y����G��X	��*���!�'�'�&�-�u��������^��1��*��
�f�y�a�~�W�W���&����_��h��@���%�u�h�}�6��(���M�Փ� F��SN����
� �`�m�'�t�}���Y����_T��h��@���%�u�h�_�w�}�W�������l ��^�����=�;�}�8��i����Lƹ��V�
N��R���9�0�_�u�w�}�W�������T��B1�@���n�u�u�%��1�(ہ�����l��S�����:�<�
�0�#�/��������C9��[\��*���`�g�%�|�|�(�����θ�C9��h��C���%�|�n�u�w�-�!���&ƹ��lP��h�I���u�u�u�u�$�1����H����S��G]�����}�0�
�8�f���������F9��1��]���h�r�r�u�;�8�}���Y���@��R�����
� �a�f�'�f�W���	����9��Z�����m�
�f�i�w�}�W���YӖ��R
��1����g�u�=�;��/����&����]	��Q��CҊ�g�e�u�u�f�t����Y���F������!�9�f�
���1���s���C9��h��F���%�u�h�&�3�1��������AN��D�����8�
�l�3��e�(��Y�ƹ�@��R
�����;�!�9�c�f�t�}���Y���C	��h�����
�m�
�d�k�}��������E��X�����0�&�2�0��2�F���&����CT�\��N�ߊu�u�:�d�1��O߁�K���@��[�����6�:�}�;�>�3�ǘ�&����T��N�� ���2�0�}�%�4�3����H����O��N��U���%�&�
�4�#�;�(��&���F��S1�����#�6�:�}�2�4�ǭ�����C	��h��C���%�|�f�|�l�W�W����ԓ�F9��1��U��&�1�9�2�4�+����Q����T��(�����d�e�|�~�"�.����Q����\��h��G��|�n�u�u�&������ד�F9��1��U��}�
�
�
�"�h�D���Y����B��B1�G���|�_�u�u�5�;�(��&���FǻN��U���&�0�
�0��l�Gϩ�����^��1��*��
�g�e�u�w�l�^ϻ�
��ƹF�N�����b�3�
�f��n�}���Y����U��V��G��u�!�
�:�>�����ە��U��^	��]���<�;�1�4��2�����ғ�u ��q(��3����y�:�<�#�:�ǫ�
����WN�N�����a�
� �b�o�-�_��Hӂ��]��G��\��u�u�'�3��j�(��E����P��h��*��l�4�1�!�'�n�(���L�֓�O��N�����<�3�
�l��o�K�������9��h[�*��:�u�
� �b�k����s���A��h��B���%�u�h�}�:��F���&����CU��X�����;�!�9�d�f�f�W�������F9��1��U��}�8�
�l�1��F݁�JӞ����T�����d�d�n�u�w�.����	�֓�F9�� 1��U��}�8�
� �a�l�����Ƹ�C9��h��A���%�|�_�u�w�8�(���H¹��lP��h�I���u�u�u�u�'��݁�&����_��N�����&�9�!�%�g�;�(��&���F�_��U���0�_�u�u�w�}�����ѓ�F9��1��N���u�&�9�!�'�i��������U��_��G��u�!�%�g��8�(��KӉ��G��^�� ��e�%�|�_�w�}�����ד�F9��1��U��_�u�u�u�w�3�!�������F��R �����!�%�3�
�c��E��Y���O��[�����u�u�u�;� �8����&��ƹF��R����
� �m�g�'�}�J�������l �� _�����'�!�%�a��2�(���A�Г�O��N�����!�%�a�3��k�(��E����^��1��*��
�g�4�1�$�1����J����P��G\����u�0�
�8�e����M����[�N��U����;�0�
�;�����H����R��G\�����}�0�
�8�e����A����O�I�\ʰ�&�u�u�u�w�}��������9��d��Uʦ�9�!�%�c�1��N߁�J���9F�N��U���2�d�4�9�-�/����&����CT��_��]���
�8�g�
�"�e�O���Q���A��N�����u�u�u�u�'�d�(�������l��=N��U���
�8�g�
�"�d�B���Y���G��W�����g�e�-�'�6�����&����O��N�����!�%�m�3��n�(��E����^��h��L���%�u�;�u�$�8�(���&����]ǻN�����8�g�
� �n�m����D�θ�C9��h��*��e�4�1�<�9�:����H����l�N�����%�
� �g�o�-�W��[����[�������:�
�:�%�$�/���O����C9��Y�����e�u�9�0�u��}���Y����G��1��*��
�f�i�u�w�}�W�������]��[�*���=�;�}�8��l����@����V�
N��R���9�0�_�u�w�}�W����ԓ�l��h_�L�ߊu�u�0�
�:�n�(���H����CT�
N�����l�'�2�d�n�}����	����@��A_��\�ߊu�u�0�
�:�n�(���H����CT�
N�����2�
� �l�g�-�W���Y����G��1��*��`�%�|�_�w�}�����ѓ�F9��1��U��_�u�u�u�w�0�(�������9�������8�
�g�'�0�l�F���P���A�R��U���u�u�u�%��1�(ہ�����l��=N��U���
�8�m�3��n�(��E����^��1����d�u�:�u�'�>�����ד�]ǻN�����8�
� �g�a�-�W��[����[�������:�
�:�%�$�/���O����C9��Y�����d�u�9�0�u��}���Y����V��P�� ���`�%�u�h�]�}�W���Y����\��h��G������u�?�3�_�������T9��^��\��r�r�u�9�2�W�W���Y�ƭ�l��D�����e�_�u�u�#�/��������F9��1��U��_�u�u�u�w�0�(�������9�������6�%�3�
�`��E��Y���O��[�����u�u�u�%�4�3����J����9F���F؊� �b�e�%�w�`�_�������9����U���
� �b�e�'�t�}���Y���� 9��hW�*��i�u�;�"�>�3�������� S��Y
�����8�g�
� �n�h����s���G��1��*���
�g�i�u�>�3��������F����*���g�
� �l�b�-�^�ԜY�Ƹ�C9��h��A���%�u�h�}�'�>�����ד�@��Z��F���2�d�l�|�]�}�W���&�ߓ�F9��1��U��w�w�"�0�w�)���&����T��N�����:�&�
�#�d�m�W�������l�N����
� �a�e�'�}�J���[ӑ��]F��^	���
�0�
�g�f�}�W�������C9��Y����
�|�u�9�2��U�ԜY�Ƹ�C9��h��A���%�u�h�&�3�1��������AN��D�����%�6�;�!�;�l�(���Tӓ��Z��SF��*���
�g�d�|�]�}�W���&�ԓ�F9��1��U��w�w�"�0�w�8����	����F9��1��U���%�6�;�!�;�l�(��PӃ��VF�UךU���8�
�a�3��h�(��E���F��R �� ���2�0�}�g�e�;�(��&���F��D�����%�6�;�!�;�l�(��PӃ��VF�UךU���8�
�c�3��j�(��E�ƿ�W9��P�����:�}�=�3��8�ǫ�
����WN��G1�*���a�d�%�|�#������ι�@��R
��E���u�g�g�6�$����N���� W�
�����e�|�|�n�w�}����KĹ��lR��h�I���!�
�:�<��8��������VN��D�����g�g�6�&��(�C���	���O�=N��U���
�m�3�
�n��E��Y����_	��T1�����}�=�3�
�>�5�_�������R��h��A���%�|�!�
�9�8��������V�I��U���
�b�3�
�n��F��T�ƨ�D��^��\���_�u�u�8��m����Kù��Z�_�����u�&�2�0��o����H����X��^	��´�
�:�&�
�!�o�D���Y����D��d��Uʡ�%�f�
� �b�h����Dӕ��l
��^�����'� �&�2�2�u�E�������O������1�4�
�:�$�����?���l�N����
� �f�c�'�}�Jϭ�����Z��R�� �&�2�0�}�e�;�(��&���F��D�����%�6�;�!�;�l�(���P��ƹF��Z��A���
�m�
�g�k�}�F������@��R
�����f�3�
�b��o�W���������T�����d�
�`�|�2�.�W��B�����h]�����b�
�g�i�w�m�W����μ�a��[��*���`�a�%�u�w�-��������9�������w�_�u�u�:��@���&����CW�
N�����2�6�#�6�8�u����ۓ��Z��SF��*���<�;�d�3��d�(��U���l�N����
� �c�f�'�}�J�������l ��_�����:�u�%�6�9�)����H��ƹF��Z��L���
�e�
�g�k�}�F������@��R
�����3�
�m�
�e�}�W�������C9��Y����
�c�|�0�$�}�G��Y���F��Z��D���&�
� �`�g�-�W��
����\��h�����'�&�/�}�>�3�Ǫ�	����U��[��G���g�|�_�u�w�)���&����P��N�U���
�:�<�
�2�)�Ǭ�
����F��P ��]���d�6�&�
�"�k�B���P����]ǻN�����g�3�
�f��o�K�������T��A�����=�3�
�<�?�u����ۋ��l0��B1�F���|�!�
�;�2�8�_�������A��H�����d�3�
�g��l�D��Y����G	�G��\�ߊu�u�8�
�c�;�(��&���F�N�����&�2�0�}�8�o����Aʹ��F�D�����%�6�;�!�;�l�(��PӃ��VF�UךU���8�
�a�;�#�;�(��&���F��Z��A���
�c�
�g�/�/��������_��G�U���!�%�a�
�"�j�O���Y����G��X	��*���!�'�'�&�-�u��������\��T��*���c�a�%�|�b�t�L���YӒ��lR��Q��Gڊ�g�i�u�d�w�5��������l0��h��B���%�u�u�%�4�3����Lǹ����RN��W�ߊu�u�8�
�`�;�(��&���F��R	��*���f�m�%�}�d�p�FϺ�����O��N�����a�
� �m�o�-�W��[����[����G���
�m�
�g�j�<�(���
����T��G�����w�w�_�u�w�0�(�������9��R��]���2�d�4�9�8�8�(݁�&�ѓ�V��[����4�
�:�&��+�(���s���G��_�� ��f�%�u�h��0�(�������_��X�����3�:�
� �n�i����s���G��]�� ��m�%�u�h�>�8�(�������l��\��U���:�;�:�e�l�}�WϪ�	����U��_��D��u�4�
�
�"�i�D���Q���W��X����n�u�u�!�'�h�(���M�ד�F�(��G���
�a�
�f�f�}�������9F���*���3�
�e�
�f�a�W���&�ޓ�F9��1��]��x�d�1�"�#�}�^�ԜY�Ƹ�C9��h��@���%�u�h�8�9�����K������^ ����� �&�2�0��0�(�������U��^��D���1�"�!�u�8�4����ۓ��Z��SF����
�4�!�3��n�(��P�ƻ�V�C�����0�}�;�<�9�9����M¹��@��B1�E���|�k�u�u�9�}����������^	��¡�%�a�
�4�#�;�(��&���[��N�����x�n�u�u�#�-�Bׁ�����l��S��G���
�a�
�g�f�}�������9F���*���3�
�m�
�f�a�W���&�Փ�F9��1��]���u�u�:�;�8�m�L���YӒ��lP��Q��LҊ�f�i�u�u�w�}�WϿ�&����G9��1�U���;�}�8�
�c�;�(��&���F�_��U���0�_�u�u�w�}�(�������9��d��Uʡ�%�c�
� �b�d����Dӕ��l
��^�����'�'�&�/��3����ے��lP��E��D��|�`�|�n�w�}����O����lS��h�I���!�
�:�<��8����
����l
��CF�����0�}�%�6�9�)���&����u ��q(��3���!�
�;�0�2�u�������A���*���3�
�a�
�f�n�Z�������V�G����u�8�
�f�1��Bׁ�K�����hX�����`�
�g�-�%�<�(���
����R��q(��3������n�w�}����Oƹ��lS��h�I���
�4�g�f�1��F݁�J����W	��C��D��u�u�!�%�a����@����[��h8��G���3�
�d�
�d�l�Z������\F��d��Uʡ�%�c�
� �a�h����DӖ��R
��1��*��
�g�f�u�8�3���P���F��G1�*���b�g�%�u�j�-�ށ�����l��_�����:�d�|�_�w�}����H����S��G]��Hʥ�&�
� �c�n�-�_������\F��UךU���8�
� �c�f�-�W��Q����S��B1�D���u�;�u�0��0�O���&����CT�=N��U���
�
� �f�c�-�W��
����\��h�����'�&�/�}�9�4��������^��h��F���%�|�d�|�l�}�Wϫ�&����F��1������3�
�e�a�-�W��s���F�G1��؊�
� �
� �n�k�������@��C��G���
�e�e�%��t�J���^�Ʃ�@�N��U���&�9�!�%�g�;�(��&����F�B"��&����!��7�%�>�(�������R��N�U���
�:�<�
�2�)�ǫ�
����WN��h�:���f�
�:�4�����HŹ��F�B �����}�;��'�8��^��Y����]��Q��*���l�a�%�u�j�W�W���Y�Ƹ�C9��h��L���%�u�=�;��8�(���Kʹ��l_��h�E���u�d�|�0�$�}�W���Y����V
��Z�*���l�`�%�n�w�}��������l��h��L���%�u�h�}�9�8����&����R��N��ʴ�
�:�&�
�!��^����Ʈ�[��=