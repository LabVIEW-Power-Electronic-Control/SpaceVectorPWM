-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǶd�����,�<�0�n�]�.�W���ݕ��l
��^��D��4�9�u� �2�4��������T��B �����{�9�n�_�9�4�ϳ�I����uV��1��*ڊ�a�
�
�
�6�}��ԜY�ƫ�]��TFךU���u�u�u�u�2�����Y����@��Y	��H���9�6�w�u�w�}�W���Y����D��_N��U��<�!�2�'�m�}�F���Y���F�N�����=�u�u�o�>�)����C����l�N��U���u�8�8�&�-�}�W������V�
N�U���|�u�u�u�'�/�W�ԜY���F�V
��E���u�o�<�u�#�����&����\��@����1�"�!�u�~�}�W���Y�����N��U���u�;�&�1�;�:����Y���F��U���u�u�u� �w�)�(�������P��
�����d�1�"�!�w�t�}���Y���F��S�U���o�<�u�!��2����������S��Dʱ�"�!�u�|�w�}�W���Y����VW�N��U���;�&�1�9�0�>�W���Y���F��N��U���u�u�;�&�3�1��������AN��^
��X���:�;�:�e�l�W�W���Y���D��N��U��<�u�!�
�8�4�L�ԜY���F�F_��U���u�o�:�!�$�9��������G	��S�����u�:�;�:�g�f�W���Y�����N��U���o�<�u�!��2����Y���F��Y
�����,�u�_�4�4�4�����ƾ�_F����L���3�e�9���Cځ�&ù��^F��d�����9�4�1�e�#�-�Mϭ�����Z��R��´�<�!�x�u�8�3���B���T����ۊ�8�u�u�!��2����������S��Dʱ�"�!�u�|�w�)��������A��^�����u�e�!�u�2�����H�ƣ���h�����0�!�'�}� �9�������\F��N�����1�#�'�4�;�}����Y����R��NUװ���<� �0�&�9�/��������@��Y	����'�7�!�u�.����� ����UF��ZN����4�9�u�&�u�1��������R��^��ʧ�8�&�,�0�m�.����B����A��C�����!�9�u�3�%�0�MϨ�����VF����*���0�_�!�'�5�)�W���0����}2��r)��!�������m�.����B���T��=d�����,�4�6�&��(����CӖ��P��F����u�7�2�;�w�}�WϿ��֓�^�
N����_�x�,�!�2�4�W�������V9��Qd��U���<�u�����2���Q����O���*���0�d�u�=�9�}�W���Y���R��1����u�:�=�'�w�c�P���B���F��[�����u�u�u�u�6�9�G���	���R��UךU���u�;�u�3�]�p��������G��D�����_�;�u�'�4�.�L���&����A��T����u�'�6�&�w�>����s����]FǻN�����9�r�#�;�w�3�W���Y���O��_��U���u�u�<�u�4�m�J���^�Ƹ�V�N��U���u�u�$�u�j�/�ǝ�7����g#��eF�����!�%�|�u�w�}�W�������U]ǻN�����3�_�;�u�%�>���s����A��T�����4�1�d�u�%�>��������F��R	�����u�u�1�'��0�W������l�D�����&�!�4�&�6�8����Y�����-��#������4�3�l�W�������I�N���ߊu�u�u�u�w�<�������F��C����u�e�|�_�w�}�W������F�N��U���'�
�8�u�j�<���s���F��SN��N���&�;�=�&�$�)��������]l��SN�����&�_�%�8�:�/�(�������	F��X�����9�|�u�7�0�3�}���Y���P
��R��ʴ�1�6�>�h�p�z�W������F���]���u�u�d�|�#�8�W���Y���F���]���u�u�d�|�#�8�W���Y���F�N��U���}������%ǿ��ד�^�T����_�u�u�u�w�}�W���Y����F�N��U���$�u�h�'�:��9���7����aN��S�����|�u�u�u�w�}������ƹF��Y
�����;�u�'�6�$�f�}��Ӕ��lǑ{�������n� �2��2�������T��_�[���n�_�;�<�.�0�G��L�֪�9��h^��Aߊ�
�u�&�u�w�:������ƹF�N�����<�!�u�u���2���D����9F�N��U���'�&��;�2�g�>���>���F��=N��U���u�1�'�&� �9���0����v4�
N�N���u�%�'�u�]�}�W���Y����GF��~ ��!�����n�u�w�}�WϽ�����}F��s1��2���_�u�u�u�w�9����I����}F��s1��2������}�3�/�������W��x9��:��n�u�u�u�w�>�G��0�Ɵ�w9��p'�����u�u�u�e�m��#ύ�=����z%��r-��'�!��1�=�z�l�3���-����l�N��Uʴ�1�0�&�u�w��$���5����l0��c!��4���0�&�<�!�w�}�W���7���]ǻN��U���0�u�u����;���:���F�N��D���u��
���L���Y�����N��U���
���
��	�%ǚ�����G�_��:����e�n�u�w�}�Wϯ�Y�ƃ�gF��s1��2������}�6�<����Y����w)��c!��\��0�1�0�!�#�f�}�������G����ʺ�u��l�g��;�G���&ù��9��N�����u�:�%�;�9�}�6��KƠ��lV��C1��A���0�e�'�8�>�W�W���Y�Ƽ�A�=N��U���u�u�u�9�w�}�9ύ�=����z%��N��U���u�u�4�1�g�g�>���-����t/��a+��:��u�u�u�u�w�}���Cӯ��`2��{!��6�ߊu�u�u�u�w�}�G��6����g"��x)��*�����_�u�w�}�W���Y����F��~ ��!�����
����}���Y���F�T�Oʜ�u��
���f�W���Y���F��N�<����
�����#���s���F�N����o��u����>��Y���F�N��D��������4���:����l�N��ʶ�8�:�0�!�]�W���������Y�3ڳ�e�9�
�
�c��(߁�����	F��X�����u��l�g��;�G���&ù��9��1�����u�%�'�u�6�}�}���Y���P
��
P�����u�u�u�u�6�9�G��Y����V��d��U���u�6�e�h�w�8�[���Y�����
P��E�ߊu�u�u�u�3�/�W�������@��=N��U���u�0�u�k�4�l�}���Y���WW�	N��Y���u�u�u�"�f�`�W���U���F��H���d�n�_�;�w�/��������lǑ