-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�l�d�d�a���(���
����GF�N�����9�u�u����;���:���F��h��U���������}���Y����G��T��;ʆ�����]�}�W�������	F��cN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�%�<���6����g"��x)��N���u�<�
�9�?��(���Y����g"��x)��*�����}�d�3�*����P���F��h��*؊�u�u�����0���/����aF�N�����u�|�_�u�w�3����&ù��	F��=��*����
����u�FϺ�����O��N�����0� �;�e�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����V��Y1�Oʚ�������!���6���F��@ ��U���_�u�u�%�%�)����Y�ƃ�gF��s1��2������u�d�}�������9F������'�
�u�u��}�#���6����e#��x<��Bʱ�"�!�u�|�]�}�W�������z(��c*��:���u�n�0�1�]�W��������A��R��U���8�l�d�d�c��(���Y���F�T�����u�%�6�;�#�1����H����g"��x)��U��r�r�_�u�w�2����Ӈ��P	��C1�����e�o�����4��Y���9F������!�4�
��$�l����I����g"��x)��*�����}�u�8�3���Y���V��L�U���6�;�!�;�w�-�$�������^9��N��1��������}�CϺ�����O�
N��E��w�_�u�u�8�.��������l��h��*���u��
����2���+����W	��C��\��u�e�d�e�l�}�WϽ�����GF��h=�����3�8�f�o���;���:����g)��Z�����:�e�u�h�u�l�G���s���P	��C��U����
�!�
�$��W���-����t/��a+��:���a�1�"�!�w�t�M���H����]ǻN�����4�!�4�
�8�.�(���K���5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��2����¹��	F��s1��2������u�g�9� ���Y���F�UךU���:�&�4�!�6�����&����lW�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��_�����u�:�&�4�#�<�(���
���� T��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��h]��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�D���_�u�u�:�$�<�Ͽ�&����G9��Y��L��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�e�d�g�l�F��H����F�T�����u�%�6�;�#�1�D݁�<����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����4�!�4�
�8�.�(���K���5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����W�=N��U���&�4�!�4��2�����ԓ�\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����W��UךU���:�&�4�!�6�����&����lV�=��*����
����u�DϺ�����O�
N��E��e�e�e�e�g�f�W�������R��V�����
�#�g�d�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�f�l�U�ԜY�Ư�]��Y�����;�!�9�f���1���?����g"��x)��*�����}�d�3�*����P���V��_�D��d�d�d�d�f�l�F��H����]ǻN�����4�!�4�
�8�.�(���K����V��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��u�u�6�;�#�3�W�������l
��1�Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[�*��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D������o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�d�d�n�w�}��������R��X ��*���g�d�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�d�e�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�d�g��}���Y����G�������!�9�d�
�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��UךU���:�&�4�!�6�����&����lW��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}��������EU��+��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��_�D���_�u�u�:�$�<�Ͽ�&����G9��1�Oʆ�������8���Kӂ��]��G��H���d�w�_�u�w�2����Ӈ��P	��C1��A���o������!���6�����Y��E���h�w�d�d�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�g�m�U�ԜY�Ư�]��Y�����;�!�9�g�g�g�$���5����l0��c!��]���:�;�:�e�w�`�U��B�����D��ʴ�
�:�&�
�!��W���-����t/��a+��:���g�1�"�!�w�t�M���H���9F������!�4�
�:�$��܁�Y�Ɵ�w9��p'��#����u�g�1� �)�W���C���V�=N��U���&�4�!�4��2�����Г�u ��N��1��������}�F�������V�S��E��d�d�d�d�f�l�U�ԜY�Ư�]��Y�����;�!�9�d��m�G��*����|!��h8��!���}�`�1�"�#�}�^��Y����V��^�E��e�n�u�u�4�3����Y����\��h��F��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I��ƹF��X �����4�
�:�&��+�(���Y����)��t1��6���u�g�1�"�#�}�^��Y����]ǻN�����4�!�4�
�8�.�(���&����`2��{!��6�����u�g�3�*����P���V��UךU���:�&�4�!�6�����&����F��d:��9�������w�o��������\�^�W�ߊu�u�:�&�6�)��������_��N�&���������W������\F��T��W��w�_�u�u�8�.��������]��[�*��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D��ي�u�u��
���(���-���F��@ ��U���o�u�e�e�l�}�WϽ�����GF��h�����#�d�f����W���-����t/��a+��:���f�u�:�;�8�m�W��[����W��_�D��d�d�d�d�f�l�F��B�����D��ʴ�
�:�&�
�!�l�C��I����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��2�����ԓ�F��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-��������lU�=��*����
����u�W������F��L�W�ߊu�u�:�&�6�)��������_��hZ��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�:�$�<�Ͽ�&����G9��1�Oʆ�������8���Jӂ��]��G��H���e�d�n�u�w�>�����ƭ�l��D�����e�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��Y����
�e�e�e�g�g�$���5����l0��c!��]��1�"�!�u�~�g�W��H����V��^�E��e�e�e�e�g�m�U�ԶY����Z��[N��*���3�8�o����0���/����aF�
�����e�u�h�w�g�m�U�ԜY�ƭ�G��B�����0�6�1�;�w�}�������F��C�� ���3�8�0�6�3�3�W�������l ��T�����9�<�u�;�9��}���Y����R
��G1�����0�
��&�f�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������	F��x"��;�ߊu�u�<�;�;�.��������lW��N�&���������W������\F��d��Uʦ�2�4�u�
�6�o�E���&����CT�=��*����
����u�FϺ�����O��N�����4�u�
�4�e�o����H����	F��s1��2������u�d�}�������9F������;�"�<�;�>����H����	F��s1��2������u�g�9� ���Y����F�D�����0�&�2�7�#�/���H����`2��{!��6�����u�e�3�*����P���F��P ��U���
�
� �g�n�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��*���
�m�b�o���;���:����g)��^�����:�e�n�u�w�.����Y����Z��D��&���!�
�&�
�w�}�#���6����9F������4�
�<�
�3��O��;����r(��N�����4�u�8�
��8�(��A����g"��x)��*�����}�u�8�3���B�����Y��������!�f�d�!�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�-������&����e9��E��D��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&�Փ�V��Z�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�;����I����	F��s1��2������u�g�9� ���Y����F�D�����9�
�0�
�o�h�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�����0�8�a�`��;�(��&���5��h"��<������}�e�9� ���Y����F�D�����-�
�:�0�#�/�(��&����T9��^��U���
���
��	�%���Kӂ��]��G�U���&�2�4�u�/��2�������9��Q��Eڊ�g�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�	����K)��h_�*���0�
�m�m�m��3���>����v%��eN��Gʱ�"�!�u�|�]�}�W�������Z��^��*���
�m�m�o���;���:����g)��^�����:�e�n�u�w�.����Y���� ^��R	��M��o������!���6�����Y��E��u�u�&�2�6�}�(���K����U�� Z��G��������4���Y����W	��C��\�ߊu�u�<�;�;�-�!���&�Փ�V��Y�Oʆ�������8���H�ƨ�D��^����u�<�;�9�9�*��������U��^��F��������4���Y����\��XN�N���u�&�2�4�w�8��������l��h_�@��������4���Y����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_�������V�=N��U���;�9�!�%�f�����A���5��h"��<������}�w�2����I��ƹF��^	��ʇ�;�0�
�9��3����&����CT�=��*����
����u�W������]ǻN�����9��;�0��1�(���
����lW��N�&���������W������\F��d��Uʦ�2�4�u�4�0�l��������l ��]�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�����&����I��D1����e�u�u����>���<����N��S�����|�_�u�u�>�3�Ϯ�M¹��U��X��G��������4���Y����\��XN�N���u�&�2�4�w��F�������
V��N��1��������}�GϺ�����O��N�����4�u�8�
��(�A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�
�0�
�n�n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h��*���$��
�!��.�(���Y����)��tUךU���<�;�9�4��4�(���&���$��{+��N���u�&�2�4�w�(�(������� 9��^�����2�
� �d�g��D��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��X��&���:�
�f�"�>�8��������T9��^��U���
���
��	�%���Y����G	�UךU���<�;�9�'��;�(��N����	F��s1��2������u�d�}�������9F������'��'�2�f�o�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��E1��G���
�e�d�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����A9��1����f�u�u����>���<����N��
�����e�n�u�u�$�:����&����lT��Q��E���%�u�u����>���<����N��
�����e�n�u�u�$�:����&����lT��E��D��u�u��
���(���-��� U��X����n�u�u�&�0�<�W�������lT��Q��E���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϱ�&����9��h��*��d�o�����4���:����V��X����n�u�u�&�0�<�W���&����l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}�����ޓ�V��Z�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)��������
S��N��1��������}�GϺ�����O��N�����4�u�0�
�:�l�(���H����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�n����H����	F��s1��2������u�g�9� ���Y����F�D�����8�
�f�3��o�@���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����g�
�0�
�n�d�Mύ�=����z%��r-��'���e�1�"�!�w�t�}���Y����R
��G1�����0�
��&�c�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������V9��E�� ���`�
�
�
�"�l�Oف�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�!��&��)��������l0��h��*��a�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�/����@9��h_�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������U��[��G��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����W��N�&���������W��Y����G	�UךU���<�;�9�!�'�n�(���H�ד� F��d:��9�������w�m��������l�N�����u�
� �d�b�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h��*���d�l�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӗ��G9��h_�*��o������!���6�����Y��E��u�u�&�2�6�}����
����9��h\�*��o������!���6�����Y��E��u�u�&�2�6�}�(���K�ד�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(ہ�����l��N��1��������}�D�������V�=N��U���;�9�!�%�1��C܁�K����g"��x)��*�����}�u�8�3���B�����Y��������!�f�j�!���&����CT�=��*����
����u�FϺ�����O��N�����4�u�4�'��(�E���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�
� �g�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h ��*��� �g�f�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������A��P��*���g�m�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӂ��V��h�����
�b�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ʈ�^��RZ�����'�4�
�
�"�o�N���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����'�
� �g�n�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E����
�
� �f�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Y
�����
� �f�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W�������	��E�����
�l�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƣ�T9��T1�����
�g�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�CW��B1�M���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l��B1�C���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'��݁�&����U��^��F��������4���Y����W	��C��\�ߊu�u�<�;�;�-�!���&ǹ��lU��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�#�-�E���&����CT�=��*����
����u�W������]ǻN�����9�3�%������@����F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�-�!�������@��h��G���%�u�u����>���<����N��
�����e�n�u�u�$�:��������`��C1�L���d�3�
�m��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��Z��B���
�f�
�d�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������^��1��*���
�f�o����0���/����aF�
�����e�n�u�u�$�:����&¹��lR��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u���F���&����CT�=��*����
����u�W������]ǻN�����9�$�<�
��(�C���	����`2��{!��6�����u�e�3�*����P���F��P ��U���4�&�2�
��(�C���	����`2��{!��6�����u�e�3�*����P���F��P ��U���4�g�d�
�"�i�C���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����d�
� �a�g�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��G1�����
�
� �`�e�-�W���-����t/��a+��:���g�1�"�!�w�t�}���Y����R
��h<�� ���`�3�
�d��i�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���a�a�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӵ��T��V�����
� �`�g�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h_�����a�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����l��N!��*��
� �`�g�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������[1��0ښ�!�d�e�3��h�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N������e� �
�b����K����	F��s1��2������u�g�9� ���Y����F�D�����8�
�a�3��j�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����1�
�0�8�d�i�!���&����CW�=��*����
����u�EϺ�����O��N�����4�u�8�
��(�B���	����`2��{!��6�����u�g�3�*����P���F��P ��U���'�
�
� �a�i����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��
�����
�0�:�
�"�k�O���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V��*���
�d�3�
�c��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��U�����<�
� �c�f�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��F���
�`�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƨ�_��S1�����
� �c�a�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������1�����a�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����A��1�����4�
�d�3��k�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
�0�:�2�9�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�
� �c�o�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Y
�����
�
� �c�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��A�����d�3�
�c��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G]�� ��`�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������T��h�����m�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����A ��@1�����3�
�e�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����C9��[\��B݊� �
� �b�`�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��G1��؊�
�c�3�
�f��D��*����|!��h8��!���}�`�1�"�#�}�^�ԜY�ƿ�T����*���3�
�g�
�d�g�$���5����l0��c!��]���1�"�!�u�~�W�W������� ��h �����'�
�`�
��(�@���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʼ�8�
� �`�b�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R�� ��e�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��Q��Aۊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���	����l �� [�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)��������9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�(���N�ӓ�F��d:��9�������w�m��������l�N�����u�0�
�8�a�9��������lQ��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����A��h��B���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	�Փ�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1�������� 9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�E�������]9��hY�*��o������!���6�����Y��E��u�u�&�2�6�}�����ғ�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����&����Q��N�&���������W������\F��d��Uʦ�2�4�u�0��0�D���&����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'����H����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�g�1��C؁�K����g"��x)��*�����}�u�8�3���B�����Y�����:�1�3�
�f��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��Y����� �m�f�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����]��R�����g�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӊ��P	��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������WT��B1�D���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1�����Փ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�8�$���&���� Q��N�&���������W��Y����G	�UךU���<�;�9�3�'��0�������l0��B1�A���u�u��
���(���-��� T��X����n�u�u�&�0�<�W���*����U��[��F��������4���Y����W	��C��\�ߊu�u�<�;�;�3� ���O����Q��G]��U���
���
��	�%���Kӂ��]��G�U���&�2�4�u�2��ׁ�����l��N��1��������}�D�������V�=N��U���;�9�;�"�2�j����Nʹ��\��c*��:���
�����o��������l�N�����u�-�
�:�2�)����L˹��P��h��B���%�u�u����>���<����N��
�����e�n�u�u�$�:��������9��hW�*��o������!���6���F��@ ��U���_�u�u�<�9�1�����ߓ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�8�$���IĹ��@��B1�B���u�u��
���(���-��� T��X����n�u�u�&�0�<�W���*����l ��\�����u��
����2���+������Y��E��u�u�&�2�6�}��������P��h��L���%�u�u����>���<����N��
�����e�n�u�u�$�:��������W��B1�M���u�u��
���(���-��� T��X����n�u�u�&�0�<�W���*����l ��[�����u��
����2���+������Y��E��u�u�&�2�6�}�����ԓ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�8�$���K¹��@��V�����c�
�f�o���;���:����g)��\�����:�e�n�u�w�.����Y����V
��h��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϰ�����9��hW�*��o������!���6�����Y��E��u�u�&�2�6�}�����ӓ�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'��݁�&����W��N�&���������W��Y����G	�UךU���<�;�9�%��1�(ہ�N����
T��G]��U���
���
��	�%���Kӂ��]��G�U���&�2�4�u�:��B���&����l��N��1��������}�D�������V�=N��U���;�9�!�%�f����H����\��c*��:���
�����n��������l�N�����u�
�4�g�d�;�(��&���5��h"��<������}�e�9� ���Y����F�D�����
�4�g�g��(�O���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʡ�%�d�
� �f�o�(��Cӵ��l*��~-��0����}�f�1� �)�W���s���@��V�����m�3�
�e�`�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��C��Dӊ� �d�f�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h[�����e�b�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӏ��CW��B1�@ߊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���	�ӓ�\��B1�Bي�g�o�����4���:����V��X����n�u�u�&�0�<�W���&�ޓ�F9��Y��G��������4���Y����\��XN�N���u�&�2�4�w�8�(���@����V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����N����\��Y1��*��d�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CW��h
�����;�3�
�d�n�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����
� �d�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���d�g�
�d�m��3���>����v%��eN��Aʱ�"�!�u�|�]�}�W�������^��1��*��e�%�u�u���8���&����|4�Z�����:�e�n�u�w�.����Y����_T��1��*��f�%�u�u���8���&����|4�Z�����:�e�n�u�w�.����Y����@��hY�� ��`�
�a�o���;���:����g)��\�����:�e�n�u�w�.����Y����Z��^��*���d�a�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƽ�]	��^\�� ��c�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����T9��h_�L���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������9��h_�D���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����K����lW�� 1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'�3��������W��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2�.�����֓�\��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������VU��^1��*��d�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������U
��h\�� ��e�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����U
��h\�� ��m�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����A ��@1�����3�
�g�l�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������R��*���g�3�
�g�d�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��A���
�g�d�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����Q��E	��*���d�g�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������9��h_�L���u�u��
���(���-��� V��X����n�u�u�&�0�<�W���&�ѓ�R��Q��G���%�u�u����>���<����N��
�����e�n�u�u�$�:����&����lU��Q��G���%�u�u����>���<����N��
�����e�n�u�u�$�:��������U��W�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�3� ������� 9��h_�C���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������U��^�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�4����H����T��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�%�8����J����U��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��C���&����l��N��1��������}�GϺ�����O��N�����4�u�
�:�d��F���&����l��N��1��������}�GϺ�����O��N�����4�u�0�&�0�?��������9��h_�M���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l��Q��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϫ�����\��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������\��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������_	��1�����
�f�m�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������A��P��*���3�
�f�g�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������V��Fފ� �d�m�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������R��F���
�f�a�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������l0��1�C���-�3�
�f�g�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1��؊�
�m�3�
�d�e����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*���
�&�$���)�(���&����`2��{!��6�ߊu�u�<�;�;�<�(���&����P��N��:����_�u�u�>�3�Ϫ�	����P��h��D��
�d�o����0���/����aF�N�����u�|�_�u�w�4����	����9��h��D��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������9��h_�M���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������G9��Q��A���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϯ�����9��h_�M���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1�����ԓ�F9��V��F��������4���Y����\��XN�N���u�&�2�4�w�/����&�ғ�F9��Z��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������V��N�&���������W������\F��d��Uʦ�2�4�u�
�8�n�(�������^��N�&���������W������\F��d��Uʦ�2�4�u�0�$�:����I����l��Q��A���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϼ����� _��1��*��a�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������U
��hZ�� ��m�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����U
��hZ�� ��`�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����A ��@1�����3�
�a�g�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������R��*���a�3�
�a�a�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h8��G��
� �d�d��l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�����3�
�a�m�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������V��D���8�-�3�
�b�i����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��#���
�
�l�3��h�E���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����6�
�4�0��/��������e9��Q��@���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l%��R1����� �0�a�
�����@Ĺ��\��c*��:���
�����l��������l�N�����u�-�
�����������G9��1�����
�`�m�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����U��T������'�6� �2�i�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�-��)�4���&����P��R1�*���
� �d�`��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��O�����&�
�!� �#�/�(���/�ғ�F9��_��F��������4���Y����W	��C��\�ߊu�u�<�;�;�;����&����l5��B�����l��m�3��h�@���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����9�
�d�
�/��$���6����F��Q��@���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l%��R1����� �0�a�
��(�F��&���5��h"��<������}�f�9� ���Y����F�D�����-�
�!��$���������T��h_�� ��m�
�f�o���;���:����g)��]����!�u�|�_�w�}����Ӏ��l��t��*��� �!�'�
�e��E���&����l��N��1��������}�D�������V�=N��U���;�9�3�%�4�����*����G��hZ��#���3�
�`�b�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��a��*��
�4�g�&�1��B���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�%�6�
�4�2���������9��Q��C���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l%��R1����� �0�`�
�����Hǹ��\��c*��:���
�����l��������l�N�����u�-�
�!��.�(�������V9��h8��*���d�g�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������K��C1�����!� �!�'��k�!�������^��N�&���������W��Y����G	�UךU���<�;�9�!�'�h�(���H����CR�=��*����
����u�W������]ǻN�����9�!�%�`��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�`�
� �f�j�(��Cӵ��l*��~-��0����}�e�1� �)�W���s���@��V�����
� �d�a��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��\�*ڊ�m�m�a�3��k�D���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����
�;�
�
�%�)�(�������F9�� _��F��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����^��GZ��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�k�(���H����CU�=��*����
����u�W������]ǻN�����9�!�%�`��(�F��&���5��h"��<������}�g�9� ���Y����F�D�����6�%�
� �f�d�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��E��
�
�m�m�c�;�(��N����	F��s1��2������u�d�}�������9F������&�1�
�;������&����T��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������9��h_�B���u�u��
���(���-��� F��@ ��U���_�u�u�<�9�1����O����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Bف�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�6�'����JĹ��\��c*��:���
�����}�������9F������%�e�b�
��e�A�������W��N�&���������W��Y����G	�UךU���<�;�9�&�3�����&����V9��D��*؊� �d�`�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������Z1�����"�<�0�4�$�:�(�������Q��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�$�9�(���&����Z��V�����
�4�!�3��j�D���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����
�;�
�
�%�)�(�������l��C1��*��l�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����V
��1����� �d�l�
�f�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����R��d1����������4���Y����\��XN�N�ߠ7�2�;�_�]�}�W��Y����P��R �����0�}�%���.�^ϱ�Y����@��RN�����0�u�x�u�w�<�(�������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N�����
�&�u�h�6��#���H����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�&�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����2�u�'�6�$�s�Z�ԜY�Ƽ�\��DN�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D����F��R ךU���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������O�C�����u�u�u�u�w�}�W����ד�_
��Y�����d�l�u�h��3�ށ�����V��B1�M���n�u�u�u�w�}�W���YӴ��T��V�����&�'�2�d�g�}�Jό�����R
��M�����
�f�
�g�]�}�W���Y���F�Q��4����!�d�l��n����H����[��O��7��� �
�c�
�����M����9F�N��U���u�u�u�-������&����e9��P1�@���h�3�%������L����F9��1��N���u�u�u�u�w�}�Wϸ�	����V9��E��Eߊ�
�0�
�m�g�a�W���&����l��Z1�@���3�
�l�
�f�W�W���Y���F�N�����;�<�
�
�2��O��E�Ƽ�e��h\�����b�
�g�d�w�2����H����F�N��U���u�u�%�a������@���F��_��*���`�c�%�n�w�}�W���Y���F��h8��G��
�0�
�m�n�a�W����ԓ� 9��hZ�*��_�u�u�u�w�}�W���Y����Q��1����c�u�h�3�'��0�������l0��B1�E���}�g�1�"�#�}�E��Y���F�N��U���8�
�d�'�0�l�N���DӒ��lW��Q��MҊ�g�_�u�u�w�}�W���Y�Ƹ�C9��h��*��e�i�u�-������&����e9��Q��@ފ�f�f�u�:�9�2�D���s���F�N��U���!�%�f�
�2��O��E�ƪ�C9��p����`��3�
�g��E��Y����G	�G�U���u�u�u�u�w�}����L����lW��N�U���4�%�4�d��n�W������O��N��U���u�u�u�u�"�)����H����[��[�� ��e�%�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�&�<�;�'�2����Y��ƹF��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����U��G��U���;�u�u�u�w�}�W���YӀ��l��t��*��� �!�'�
�a��@�������F���*����&�
�!�"�)����O����l ��]�*��_�u�u�u�w�}�W���Y����U��R	��L��i�u�8�
�d�;�(��N����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�}�W��Y����T��E�����x�_�u�u�%�>��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�r�p�}����Y���F�N�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����d�h�4�
�2�}��������C9��V��Hʴ�
�:�&�
�8�4�(���P�Ƹ�VǻN��U���u�u�u�u�2�.��������lW��N�U���4�g�g�3��l�(��J�ƨ�D��]�N���u�u�u�u�w�}�WϮ�/����9��P1�E���h�%��9�����L����9F�N��U���u�u�u�<�9�4�(���&����Z�G1��؊�
� �d�`�'�u�AϺ�����P�=N��U���u�u�u�u�w�0�(ف�����Q�
N�����3�
�g�
�e�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߊu�u�x�4�$�:�W�������K��N�����0�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��D���!�0�_�u�w�}�W���Y���N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��h��*���|�!�0�_�w�}�W���Y���F��h��ۊ�e�'�2�d�c�}�Jϱ�&����9��h��D��
�g�_�u�w�}�W���Y���\��d�����f�"�<�0�6�.��������V�
N�����6�:�
�f� �4����
����U��^����u�u�u�u�w�}�W���	����9��h��*��c�i�u�
�6�o�Eׁ�����9��d��U���u�u�u�u�w�/�!�������
U��S��*���
� �d�f��o�}���Y���F�N�����'�2�d�g�w�`��������Q��UךU���u�u�u�u�w�}��������A��W�U��&�9�!�%�f�;�(��J����9F�N��U���u�u�u�0��0�F܁�����T�
N�����%�f�3�
�f�l���Y���F�N��U���0�
�8�m�%�:�F��Y����V
��Z�����e�`�%�n�w�}�W���Y���F��Z��*���
�l�f�i�w�0�(ׁ�����l��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}���Y���G��Y��U���!�u�4�
��;����Ӓ����C�����;�{�x�_�w�}����&����R��P �����o�%�:�0�$�u�������R��d1�����%�6�|�u�w�?����Y���F��V������3�8�<�]�}�W���Y���D����&���!�
�&�
�w�c�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�4�
�#�/�W���	����@��X	��*���|�u�=�;�w�}�W���Y���F�N�����
�&�u�h�6��#���K����lW��N��U���u�u�u�u�2�.�}���Y���F�N��U���4�
��3�:�a�W���*����9��Z1����u�u�u�u�w�}�W���Y����F�N��U���"�0�u�%���݁�
����X�N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���%��
�&�w�`����-����l ��h\�U���u�u�u�u�w�}����s���F�N��U���u�u�4�
��;���Y����g9��1����_�u�u�u�w�}�W���Y����Z ��N��U���u�u�"�0�w�-�$�������^9��
P��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}�W�������F�N��U���u�u�u�u�6��$������R��c1��F���8�g�_�u�w�}�W���Y���V��^�U���u�u�u�u� �8�W���*����9��Z1�H���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W���Y����_��N��U���u�u�u�u�w�}����*����Z�V��!���a�3�8�f�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����g9��1����h�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y���F��[��U���u�u�u�u�w�}�W�������l ��R������&�`�3�:�i�}���Y���F�N�����<�n�u�u�w�}�W�������\��E��K���u�u�u�u�w�}�W�������l ��R��W����w�_�u�w�}�W���Y����l�N��ʥ�:�0�&�_�w�}����H����l	��D1��*��
�g�i�u�f�}����Q����@��h[�� ���m�%�u�u�'�>�����ғ�F��D��E��u�u��;�2���������U��Z��G��u�d�u�=�9�u�(�������l ��_�����u�%�6�;�#�1�C��Y����D��d��Uʇ�;�0�
�9��3����&����CT�
N��Wʢ�0�u�%��$�1�(ׁ�����l��
N��*���&�
�#�
�~�8����I��ƓF�C�����;�u�&�<�9�-����
���9F������
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9�������4�
�<�
�$�,�$���ƹ��^9��=N��U���<�_�u�u�w�}����Q������T�����2�6�d�h�6�����P�ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�����e�|�:�u��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�h����M�����YNךU���u�u�u�u�'�9����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����:�0�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�4�
�1�2�<����Y����V��C�U���4�
�1�0�6�.���������T��]���&�4�!�u�'�.��������l��h��*���u�u�7�2�9�}�W���Yӏ��N��CF�����;�!�9�2�4�l�JϿ�&����GO�V ��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�~�}����s���F�N�����1�0�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӇ��Z��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����4�&�2�u�%�>���T���F��h�����&�<�;�%�8�}�W�������R��RB�����2�6�0�
��.�B������F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���ځ�
����O��_�����u�u�u�u�w�-���� ���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�'�4�,�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R�����u�4�
�0�"�3�G��Y����l��h8�����
�&�<�;�4�.�(���H����CW��N�����0� �;�d�k�}��������l��C�����;�d�6�&��(�F��&����F�V�����;�g�i�u�$�0����/����G��D�����6�&�
� �f�j�(��s���R��R����i�u�0��;�o�(�������U��h����u�x�u�%�$�:����H����@��YN�����&�u�x�u�w�<�(���&����T��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��D��i�u�4�
�8�.�(���&���R��d1����1�"�!�u�~�f�W�������A	��D����u�x�u�%�$�:����K�ƭ�@�������{�x�_�u�w�-�������� 9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�U��}�%��
�$�u�W������F�V�����
�#�
�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(������]F��X�����x�u�u�4��4�(���&�ޓ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��N�U´�
�:�&�
�!��W���	����U��N�����u�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�j�FϿ�
����C��R��U���u�u�4�
�>�����O¹��@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9��N�U´�
�:�&�
�!��W���	����U��N�����u�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�d�W�������A	��D�X�ߊu�u�%�&�0�?���&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����
P�
N�����;�!�9�d�f�`����*����T��X����|�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���ށ�
����R��P �����&�{�x�_�w�}��������B9��h��*���
�
�&�<�9�-����Y����V��V�����1�
�f�_�w�}����s���F�^�����<�
�1�
�d�}����s���F�N�����<�
�&�$���ށ�
����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����U��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�V�����&�$��
�#�����Y����T��E�����x�_�u�u�'�.��������l��h��*ۊ�&�<�;�%�8�}�W�������R��^	�����m�_�u�u�2�4�}���Y���Z �V�����1�
�m�u�?�3�}���Y���F�V�����&�$��
�#�����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�<�
�&�&��(���&����F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��^	������
�!�
�$��W�������A	��D�X�ߊu�u�%�&�0�>����-����l ��h\�����;�%�:�u�w�/����Q����Z��S
��C�ߊu�u�0�<�]�}�W���Y���R��^	�����c�u�=�;�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�1��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�
�&�
�w�.����	����@�CךU���%�&�2�6�2��#���M����lU��D�����:�u�u�'�4�.�_���
����W��\��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��D��u�=�;�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��F1��*���
�&�
�u�$�4�Ϯ�����F�=N��U���&�2�6�0��	��������l��^	�����u�u�'�6�$�u��������lQ��d��Uʷ�2�;�u�u�w�}��������T9��S1�D���=�;�_�u�w�}�W���Y����Z��D��&���!�
�&�
�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h��*���$��
�!��.�(���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�2����<é��lW��h��@���%�u�h�}�:��(���&�����������!�9�d�d�l�}�Wϼ�����vV��C1�E���
�`�
�g�k�}����J����T9��^�����%�6�;�!�;�l�F��Y����\	��O)��:���d�a�3�
�a��E��Yۓ��l��h_�@ʭ�'�4�
�:�$��ށ�P���F��Z��؊� �d�g�
�e�a�WǱ�����D9��Q��D���%�u�'� �3�/����K����l ��\�*��n�u�u�7�:�/����¹��lW��1��U��}�
�:�f��l����J�ғ�F�� �����7�!�e�;�#�4�(���H����CT�=N��U���0�2�f�
�e�;�(��M����[�G1�����<�
� �d�a��Eϱ�Y����Z��^��*���
�g�3�
�c�o����s���Q��E	��L���3�
�g�d�'�}�J���&����9��Q��D���%�u�'�;� �4����&ù��G9��Q��D���%�|�_�u�w�/����J����U��h�I���:�0�3�:�����K����	��B �����"�f�;�!�1��D���	����F�U�����e�1�8�'�6��F���&����CT�
N�����2�7�!�d�%�:�F��Y����W��C�����
�
� �c�c�-�^�ԜY�Ʈ�^��RZ�����'�4�
�
�"�o�N���Y���]��^	�����0�
�m�e�6�9��������]��Q��B؊�f�n�u�u�5�0����I����F9��1��U��}�'�0�2�c���������l ��W�����:�u�%�6�9�)����H��ƹF��E�����3�
�a�m�'�}�J�������\��h��D���
�g�:�u�9�8����&ǹ��G9��h_�G���|�_�u�u�%�8��������l��S�����
� �f�m�'�}�ϼ�����V��R�����<�3�
�l��o�L���Yӄ��V��h�����`�
�g�i�w�3� �������9��P1�M���'�%�;�!�>����L����l�N�����0�<�
� �f�j�(��E����V��P �����3�
�d�b�'�}�Ϯ�����9��h_�@���|�_�u�u�%�8����J����U��h�I���;�"�<�;�>��(���H����CU��EN�����<�
� �d�g��E��Y����A��P��A���
�a�a�%�w�`�_���
����Z��h��D��
�f�:�u��2�(������� ^��G�U���7�8�'�0�>�;�(��&���F��R�����!�'�2�d�f�}�Ϯ�����l ��V�����_�u�u�'�2�:�(���H����^��G\��H���;�0�3�:�����M����\��A�����d�3�
�c��o�L���Yӄ��V��h��G���
�g�f�%�w�`�_�������D9��Q��G���%�u�'�:�2�;����&����^��G\����u�'�0�2���D���&����l��S�� ���'�9�"�f�1��D���	�ƣ�	��E�����3�
�f�g�'�t�}���Y����A��^1��*���d�m�
�g�k�}��������lR��B1�Mڊ�g�:�u�#�%�1� �������P��G�U���7�8�'�0�>�4����HŹ��Z������:�
� �f�g�-�W�������_	��Q��Lي�g�n�u�u�4�/��������9��R��]���
�m�'�2�f�j�W���Y����W��R	��M��n�u�u�6�%�$����O����Z������
�0�
�b�b�<�Ϫ�	�Г�V��_�N���u�1�9�!�3�2����&���� R��N�U���u�u�u�%�c��(���&������YN�����
�
� �c�c�-�_���D����F��D��U���u�u��;�2���������V��W����u�0�0�0��3����&����CU�
NךU���u�u�8�
��(�E���	�ƻ�V�T�����
�c�
�g�g�}�W��PӃ��VFǻN��U���<�;�<�
�2��@��s���W��C�����&�3�
�g��n�K���Y���F��V ��D���9�:�0�
�2��O��������E��*���c�a�%�}�~�`�P���Y����l�N��Uʇ�;�0�
�9��8��������U��N��������!�f�j�!���&����CT�
N�����2�6�#�6�8�u��������C9��Y����
�|�x� �$�:��������[��h8��N���u�3�%������@����l ��V�����h�_�u�u�w�}����;����G9��1��F���
�`�
�f� �8�WǪ�	�ԓ�F9��1��]���h�r�r�u�;�8�}���Y���U��v,��:���d�l��3��j�(��s���U��v,��:���d�l��f�1��Bہ�J���9F�N��U���4�g�a�8�/�;�(��&����[�������
� �f�a�'�u�^��^���V
��d��U���u�%��9�����N����9F���*���-� �
�c�����O����[��C
�����
�0�!�'�"�.����Q����\��h��G��u�u�;�<�9�9����8����F��W��*ي� �f�a�%�~�f�W�������v!��B��Fߊ�
� �a�e�'�}�Jϭ�����Z��R�� �&�2�0�}�'�>��������O������1�3�%�;�3�����M�ӓ�l ��W�����n�u�u�3�'��0�������l0��B1�A���u�h�&�1�;�:��������F��P ��]���6�;�!�9�d��^������]��Q�����
�0�8�f�c�����@¹��O��N�����6�
�4�0��/��������e9��Q��@���%�u�h�_�w�}�W�������l%��R1����� �0�`�
������@����[����*���m�'�2�d�c�u�^��^���V
��d��U���u�3�%�6��<��������A��1�����`�b�%�n�w�}��������@��C�����
�g��g�1��B���	���l�N��Uʳ�%�6�
�4�2���������
9�� 1��*���e�%�u�=�9�u��������A��W�]���h�r�r�u�;�8�}���Y���U��T������'�6� �2�i�(���&����^��G]�U���u�u�3�%�4�����*����G��hZ��#���3�
�f�b�'�}�Jϭ�����Z��R��§�&�/�}�<�9�9����K����T9��W��F���n�_�u�u�/�����
����A��B��A؊�
�
� �d�n��D��Y���F���*����&�
�!�"�)����K����l ��]�*��"�0�u�&�;�)��������
P��G��U��|�0�&�u�w�}�W�������G9��D�����!�'�
�g��o����L�֓� ]ǻN�����!��&�
�#�(����&�ԓ�l ��[�*��i�u�u�u�w�}��������@��C�����
�g��b�1��D���	�ƻ�V�X�����
�e�'�2�f�i�_���D����F��D��U���u�u�%��;��F܁�����f$��B�� ���3�
�`�`�'�f�W�������G9��D�����!�'�
�l��n����L�ғ� F�d��U���u�3�%�6��<��������A��1��B���
�f�b�%�w�5��������C^��R	��L��e�u�u�d�~�8����Y���F��O�����&�
�!� �#�/�(���/����S��h����u�-�
�!��.�(�������V9��h8��*���d�c�
�f�k�}�W���Y����K��C1�����!� �!�'��k�!�������
Q��@��U¦�9�!�%�d�%�:�F��Q���A��N�����u�u�u�u�1�-��������G��C��*����f�3�
�b�i���Y����K��C1�����!� �!�'��d�!�������V��N�U���u�u�u�%��1�(��&����U��^�����=�;�}�'�2�:�C���&����l��G��U��|�0�&�u�w�}�W���	����9��W�� ��d�
�f�_�w�}��������V9��E�� ���a�
�
�
�"�l�A؁�J���9F�N��U���
�!��&��)��������l0��h��*��a�"�0�u�$�1����J����lW��F�U���d�|�0�&�w�}�W���YӀ��l��t��*��� �!�'�
�n��C���&����l��=N��U���
�!��&��)��������l0��B1�A݊�f�i�u�u�w�}�Wϸ�	����p��h=�� ���'�
�l��`�;�(��I����D��F��*���1�
�e�'�0�l�C���P���A�R��U���u�u�u�3�'�%�"�������Q��T��L܊�
�
� �d�e��D�ԜY�ƪ�C9��h-�����'�6� �0�b��(݁�����9��R�����u�u�u�-��)�4���&����P��R1�*���
� �d�g��n� ���Yە��l��1����a�}�|�h�p�z�W������F�N�����
�4�0��%�>����LŹ��U��^����u�u�3�%�4�����*����G��h[��#���3�
�c�d�'�}�J�ԜY���F��G1��*���0��'�6�"�8�C݁�&Ĺ��lW�� 1��U���;�}�0�
�:�l�(���&����V�
N��R���9�0�_�u�w�}�W���&����R��d�����0�`�
�
��(�F��&����F�Q�����4�0��'�4�(���&����U��V�����h�_�u�u�w�}�(���K����l��h��D��
�f�"�0�w�?��������lW��1��]���h�r�r�u�;�8�}���Y���C9��[\��*���3�
�f�m�'�f�W�������G9��D�����!�'�
�c��e����O�ޓ� F�d��U���u�3�%�6��<��������A��1��B���
�`�e�%�w�5��������CW��E��D��}�|�h�r�p�}����s���F�Q�����4�0��'�4�(���&����U��\����u�u�3�%�4�����*����G��h[��#���
�c�m�%�w�`�}���Y���U��T������'�6� �2�h�(���&����_�������'�6�;�d�e�����@���F�_��U���0�_�u�u�w�}�(���K����l0��1�����`�d�%�n�w�}�W�������\��C��*��
�
� �`�f�-�W��
����\��h�����'�&�/�}�>�3�Ƿ�&����R9��aG�F���_�u�u�u�w�;��������A��[��*���f�c�%�u�j�.��������V��EF�����}�<�;�1�1�-�6���6����_��h]�� ��a�%�|�f�~�f�}���Y���U��Y��*���8�a�m��4�.�(���N�ѓ�F���*���<�
�0�!�%�/����Q����V��O�����!�'�
�`�����@����U��UװU���3�%�;�1��8���A����F9��1��U��}�8�
�a�1��Eށ�J����C9��Y����
�|�_�u�w�%�(���;����l5��C����c��&�3��h�O���Y���F�N�����6�
�4�0��/��������e9��Q��@���%�u�=�;��0�(ׁ�����U�N��R��u�9�0�_�w�}�W�������l%��R1����� �0�a�
�����@Ĺ��l�N����
�:�
� �f�j�(��E����P��h��D���
�g�-�'�6�����&����O��N�����d�3�
�e�b�-�W��[����[����*���3�
�e�b�'�}�W�������l
��h^�����u�d�n�u�w�4��������_��N�U��u�=�;�}�>�3�Ǫ�	����U��]�����i�&�2�0��-��������lW������w�_�u�u�4�-�(���H����CT�
N��Wʢ�0�u�&�2�2�u����@����P��h�U���<�;�1�4��2����ǹ��F��D��E��u�u�<�8�c�;�(��N����[�L�����}�<�;�1�#�-�Aށ�����9��N����0�}�%�6�9�)����H����_��^�����u�6�%�3��e�(��E���F��R �����f�
� �`�`�-�W���	����@��A\��\ʰ�&�u�e�n�w�}����&����U��W��G��u�<�8�
�"�h�B���Y����R��X ��*���
�|�_�u�w�.����&����Q��G]��Hʥ��9�
�f�1��E���	������Y��F���_�u�u�&�2��(���H����CU�
N��#���
�d�3�
�c�n����Jӂ��]��]����u�&�0�
�"�l�Dց�J���C9��[\��E���
�d�f�%��i��������]ǻN�����'�
� �g�n�-�W��Q����Q��E��D��u�;�u�0�$�:��������W��d��Uʻ�2�&�6�;�#�;�(��&���F��R	����� �g�l�%�w�2�W�������l
��h_����u�0��9�g�;�(��&���FǻN��U���;�4�%�4�f�� ���Yە��l��1��*��
�g�e�u�w�l�^ϻ�
��ƹF�N������-� �
�a��(܁����� U��N�����0�d�
� �n�e����D���F�N�����1�
�0�8�d�i�!���&����CW��_��]���
�8�b�3��j�(��I���W����ߊu�u�u�u�/��2�������9��Q��Lފ�g�_�u�u�2���������9��R�����u�u�u�-������&����e9��h[�*��"�0�u�<�:����L����O�I�\ʰ�&�u�u�u�w�}����7����F��[��*���
�m�m�_�w�}�����Փ�F9��1��U��_�u�u�u�w�8�$���H¹��@��B1�A���u�=�;�}�%�>��������l��G��U��|�0�&�u�w�}�W�������_W��Q��FҊ�f�_�u�u�2���������9��R�����u�u�u�%�4�3����J����[����*���b�3�
�b��o�G���Y�����RNךU���u�u�%�6�9�)����K���F��@=��Dߊ� �l�`�%�w�`�}���Y���R��X ��*���
�u�=�;��>����&����CT�N��R��u�9�0�_�w�}�W���	����@��A]��N���u�;�"�0�f����J����[�N��U���;�"�0�g�f�>��������F9��1��U���;�}�'�6�9����@����O�I�\ʰ�&�u�u�u�w�}��������U�� Y��F�ߊu�u�0��;����L����[�N��U���3�%����)�F���/����lW��N�����&�9�!�%��(�@���	����[�I�����u�u�u�u�w�;��������A��[��*���
�m�e�_�w�}�W�������V��T��*���l�b�%�u�j�.��������V��EF�����}�<�;�1�9�*��������9��B�\��_�u�u�u�w�8�$���H¹��@��B1�A���u�h�&�1�;�:��������A��M�����1�;�"�0�f����A����U��UװU���;�"�0�g�f�>��������F9��1��U��_�u�u�u�w�-��������lW��_��]���
�8�`�3��m�(��I���W����ߊu�u�u�u�'�>�����Փ�l�N�����g�l�6�&��(�F��&���F��S1�����#�6�:�}�2�4�ǫ�
����WN��C1�����
�f�"�<�2�<����&����_��B�\�ߊu�u�0��;����N����[�N��U���3�%����)�F���/����lW��N�����<�8�
� �b�h����P���A�R��U���u�u�u�3�'�3��������S��h��*��e�_�u�u�2��܁�����l��S��U���u�u�;�"�2����J����D��F��*���1�3�
�d��o�G���Y�����RNךU���u�u�0��;����L����9F� ��&���
� �l�f�'�}�J�ԜY���F��G1�����0�8�a�m��>��������l��@��U¦�9�!�%�
�"�e�@���Q���A��N�����u�u�u�u�1�-�6���6����_��h]�����m�f�_�u�w�8�$���&����S��N�U���u�u�u�3�'�3��������S��h��*��e�"�0�u�$�1����&����Q��F�U���d�|�0�&�w�}�W���YӀ��l(��O!��*��
�
� �`�c�-�L���Yӈ��`��h��M���%�u�h�_�w�}�W�������t��C1�@���'�2�d�`�w�5��������CQ��B1�D���}�|�h�r�p�}����s���F�Q�����
�0�8�f�c�����@¹��l�N�����b�3�
�b��n�K���Y���F��O�����!�'�
�m�����H����D��F����� �`�`�%��t�J���^�Ʃ�@�N��U���3�%����)�F���/����_��G\�U���;�"�0�m�1��O؁�J���9F�N��U����9�
� �o�h�������\��X �����d�
�g�e�w�}�F�������9F�N��U����9�
� �o�o���Y����V��[W�� ��e�%�u�h�]�}�W���Y����V
��Q��Eي�f�"�0�u�8���������
9��^��H��r�u�9�0�]�}�W���Y����r$��x��D����f�'�2�f�n�L���Yӈ��`��Q��Dي�f�i�u�u�w�}�Wϸ�	����V9��E��Eߊ�
�0�
�m�g�*����
����^��Q��E݊�g�e�u�u�f�t����Y���F���*���-� �
�f������A����F�Y�����<�
�
�:��l����J�ޓ�F�F�����;�<�
�
�"�l�Oف�JӞ����T�����d�d�n�u�w�3� �������9��C1��*���d�c�
�g�k�}��������G9��Q��A���%�u�:�u�'�>�����ד�]ǻN�����2�7�!�e�9�)����&����l��S�����<�;�<�
��(�F��&����\��G1�����9�d�d�n�w�}��������G9��Q��Mڊ�f�i�u�
�6�o�E܁�����l��[�����:�d�|�_�w�}��������lT��B1�A݊�f�i�u�
�6�o�D߁����� 9��]����!�u�d�n�w�}��������G9��Q��G���%�u�h�%��1�(�������_��F�U���;�:�f�|�]�}�W���
����Z��h��D��
�f�i�u��<�E��&����V��G\��Dʱ�"�!�u�d�l�}�Wϰ�����Q��Q��Gۊ�f�i�u�
�6�o�E���&����CT�N�����u�d�n�u�w�2�(�������@��Y1��*���
�f�i�u�w�}�W�������C��1�����u�!�%�3��i�(��I���W����ߊu�u�u�u�/��5�������9��Q��Aӊ�g�_�u�u�%�>����Kù��lW��1��U��}�6�%�
�"�l�Bځ�KӇ����h��C���%�|�_�u�w�/����H����U��G\��H���0�
�8�b�1��@ށ�KӉ��@��C��*���b�b�%�|�]�}�W�������l ��[�����h�}�'�6�9����@����\��E1�����3�
�f�
�e�f�W�������]��B1�L���u�h�}�0��0�B���&����CT��EN�����%�
� �b�n�-�^�ԜY�ƣ�G9��T��*���"�<�0�4�$�:�(���H����CU�
NךU���u�u�0��;�k����@������YN�����;�g�3�
�b��E��Y���O��[�����u�u�u�0��1�B���&����CU��N�����3�:�
�
�"�k�F���Y���Q��E	��ۊ� �c�d�%�w�3�W���&�Փ�F9��1��\�ߊu�u�#�'�;�*�E���&����l��S�����'�0�<�
�"�l�@ށ�KӇ����h\�����d�b�%�|�]�}�W�������lU��B1�G؊�g�i�u�7�:�/����&���� W��G\�����8�
�a�3��n�A���P���F��R�����
� �d�`��o�K�������T��1��*��a�%�u�;�w�0�(�������V��G�U���:�0�3�:��(�E���	���N��Z�����3�
�m�
�e�<�Ϫ�	����F9�� 1��\�ߊu�u�
�g�d�m�G��&ǹ��lW��1��U��_�u�u�u�w�-��������9��@��U¡�%�`�
� �f�h�(��I���W����ߊu�u�u�u�:��C���&����l��=N��U���g�f�e�e�`��(���H����CU�
NךU���u�u�%�6�9�)���&�ƻ�V�C��Cڊ� �d�l�
�d�m�W���H����_��=N��U���u�8�
�`�1��A���	��ƹF��h^�F���e�m�
�
�"�l�Bށ�J���9F�N��U���6�;�!�9�d��W����θ�C9��h��D��
�f�e�u�w�l�^ϻ�
��ƹF�N�����c�3�
�c�b�-�L���YӖ��9��Q��Aڊ�g�i�u�6�%�$�F���&����CT��Y
�����d�4�9�:�2�����A���9F���D���3�
�a�
�e�a�Wǌ�����R
��X ��*���`�g�%�u�9�}����K����R��G\����u�
�0� �#�h����H˹��Z�Q��;����!�d�`��;�(��&���F��@ ��U��n�u�u�%��.����&����S��GZ��Hʥ��9�
�e�1��F���	������Y��F���_�u�u�
�2�(��������9��R��������!�f�h�!���&����CT�N�����u�e�n�u�w�-�!���&����^��Q��E݊�f�i�u�u�w�}�WϿ�&����G9��X��3���"�0�u�7�:�/����¹��lP��h�E���u�d�|�0�$�}�W���Y����l0��1�*���
�m�l�_�w�}�(���K����U��Z��A��u�-�
��/�(�(��&����lR��h�G���:�;�:�d�~�W�W���&����lW��h��*���d�b�
�f�k�}�W���Y����C9��Y����
�����*��������T��h�����f�g�%�}�~�`�P���Y����l�N��Uʥ��9�
�a�1��E���	��ƹF��h8��G��l�8�-�3��h�C���Y���F�N�����:�&�
�#�e�j�1���?�ƻ�V�U�����<�<�
� �f�e�(��I���W����ߊu�u�u�u��<�E��&����W��G_�U���%��9�
��(�F���	�����V�����
�a�
�g�c�}��������l�N��#���
�d�
�4�e�.����L�ד� F�d��U���u�3�%�6��<��������A��1��B���
�f�b�%�w�5��������A��W�]���h�r�r�u�;�8�}���Y���U��T������'�6� �2�h�(���&����_��d��Uʥ��9�
�d��%�(���;����l5��C1��*���`�%�u�h�]�}�W���Y����P��V��&���6� �0�`���(���&������YN�����
�0�
�l�d�m�W���H����_��=N��U���u�-�
�!��.�(�������V9��h8��*���d�g�
�f�]�}�W����ԓ� 9��hZ�*��i�u�!�
�8�4�(�������]��Y�����9�
�m�3��l�(��Y�ƹ�@��R
�����e�3�
�b��l�^�ԜY�Ƽ�e��h\�����`�
�f�i�w�}�W���Yӈ��`��h��M���%�u�=�;��/����K����S��G\��\��r�r�u�9�2�W�W���Y�Ƣ�D5��1��*��
�f�_�u�w�����K˹��lW��1��U��&�1�9�2�4�+����Q����V��h8�� ��d�
�g�u�w�4��������
9��h_�B���|�n�u�u�'��݁�&�ޓ�F9�� V��F��u�u�u�u�w�<�(���
���� T��^�E��"�0�u� �3�/����J����U��h�E���u�d�|�0�$�}�W���Y����l0��1�*���d�m�
�d�]�}�W����ԓ�l ��_�����h�&�1�9�0�>�����ι�@��R
��*���g�d�3�
�a��C���Y����T����*ފ� �g�d�%�~�f�W���	����9��h��D��
�g�i�u�#�����&����\��^	��¡�%�g�
� �f�o�(��Y�ƿ�T����*���3�
�d�e�'�t�L���YӖ��R
��]�� ��c�
�g�i�w�)�(�������P�������!�%�f�
�6�)����K�ӓ�O������'��'�2�f�o�^��Y����l0��1�*���d�m�
�d�k�}�(���K����U��X�����g�x�d�1� �)�W���s���C9��[\��*���3�
�`�g�'�}�J�ԜY���F��h�����#�g�m�e�g�m�W����ι�W��[��A���
�a�e�%��t�J���^�Ʃ�@�N��U���%��9�
�e�;�(��O����9F������f�3�
�l��n�K���Y���F��R��Ҋ� �m�b�%�w�5��������WT��B1�D���}�|�h�r�p�}����s���F�Y�����3�
�b�
�d�W�W���&����lR��Q��A���%�u�h�&�3�1��������AN��P ��]���
�l�6�&��(�F��&���F��P ��]���
�
�0�
�n�m�^�ԜY�Ƽ�e��hZ�����a�c�%�u�j�-�!���&�ד�F9��]��G��u�u�u�:�9�2�G��Y����l0��1��D݊� �l�d�%�w�`�}���Y���]��R�B���&�
� �l�`�-�W����Σ�l��S\�� ��d�%�}�|�j�z�P������F�N��������!�f�h�!�������]ǻN��*���g�a�3�
�c��D��Y���F������!�9�f�
�g�m�G��������R����� �f�e�%��t�J���^�Ʃ�@�N��U���%��9�
��8�(��M���F��a��*ފ� �
� �f�g�-�W��s���F�V�����
�#�g�b���1������Q��E	�����3�
�d�
�e�m�W���H����_��=N��U���u�
�4�g�e�/���I��ƹF��h8��G���3�
�c�
�d�a�W���Y�����d��F���
�`�
�f� �8�WǱ�&����9��hV�*��e�u�u�d�~�8����Y���F��R�����3�
�a�
�d�W�W���&����l��1��*��
�f�i�u�w�}�W�������]��[�*��e�"�0�u�"�9�����ד�F9��1��]���h�r�r�u�;�8�}���Y���C9��[\��F���2�d�b�n�w�}��������U��[��E��u�;�7�!���L���YӖ��R
��D1��*��
�g�i�u�#�����&����\��R�� �&�2�0�}�#�����&����\��^	��¥��9�
�
�"�l�B���P����Z��SF��R���%�6�;�!�;�i�(���N���R��UךU���
�:�f�
�f�;�(��M����[�L�����}�8�
�
�"�l�Nہ�M����C9��Y�����f�u�9�0�u��}���Y����GU��^\�� ��c�
�g�i�w�m�W����θ�C9��h��D��
�a�h�4��2����������RN��W�ߊu�u�
�:�d��(���H����CT�
N��Wʢ�0�u�%��$�1�(؁�����9��S�����;�!�9�f�`�}����[����F�G1�����
� �c�`�'�}�J�������W9��E�����g�
�f�-�%�<�(���
����9��d��Uʥ�;�!�<�
�"�l�Aځ�K���V�@��U¥��&�9�
��(�F��&�����T�����f�e�u�9�2��U�ԜY�Ƽ�]	��^]�� ��e�
�g�i�w�m�W����θ�C9��Q��G���%�u�u�%�4�3����K���V
��L�N���u�%�;�!�>����J˹��Z�^�����u�!�%�g��(�F��&�����T�����g�e�u�9�2��U�ԜY�Ƽ�]	��^1��*��
�g�i�u�$�:��������_��O�����,�3�
�c��o�L���Yӗ��R��P ��*���g�`�%�u�j�u�(���&����
_��N��ʤ�<�
� �d�d�-�^�ԜY�ƽ�l��^	��F���
�c�
�g�k�}����¹��lR��h����$�<�
�
�"�i�C���P���F��^��*���a�a�%�u�j�;����>����lW��h8�� ��e�%�}�g�3�*����K��ƹF��U�����b�
�f�i�w�����
����R��G\��Aʱ�"�!�u�a�l�}�WϬ�H����U��G\��H���w�"�0�u�#�-�D؁�����l��
N��*���&�
�#�g�g�}����[����F�E1��G���
�e�d�%�w�`��������l��C�����0�}�8�
�`�;�(��J����M��^	��¡�%�d�
� �f�o�(��P���F��a1��*��b�%�u�h�$�9��������G	��D�����8�
�`�3��m�N���P����Z��SF����
� �d�d��l�^�ԜY�ƾ�U��[��G��u�e�u�=�9�u����L����^��G_��U���6�;�!�9�f��^ϻ�
���]ǻN��*���d�3�
�`��o�K�������
9��hZ�*��:�u�
�
�"�i�A���P���F��^1�����l�
�g�i�w�)���&����
W��N��U��� �d�`�%�~�W�W�������lP��h�I���7�:�
��.�(�(��&����T��N��ʴ�
�:�&�
�!��^�ԜY�ƿ�_9��G_�����e�b�%�u�j�u��������l��X�����
�e�d�%�w�2�W�������l
��h_����u�0�
�8�f����I����Z���*ۊ� �c�c�%�w�3�W���&����9��h_�B���|�_�u�u�2����&����W��G\��H���0�
�8�d�c�9��������lW��1��U���u�%�6�;�#�1�F��B�����h��D���1�8�'�4��(�F��&���F��E1�����g�
� �d�a��Eϱ�Y����^��B1�C݊�g�n�u�u�$�1����J����\��Y1��*��
�g�i�u�$�1����&����A��h��B���%�u�'�!�'�l����IŹ��]ǻN�����8�d�
� �f�o�(��E����^��h��C���%�u�;�u�2����&����W��G\����u�0�
�8�f�i��������U��^�����h�}�0�
�:�l�@�������]9��h_�D���u�'�!�%�f�;�(��&���9F���*���d�3�
�a��o�K�������U��[��Gʭ�'�4�
�:�$��ށ�P���F��[1�����1�8�'�4��(�@���	���N��[1�����1�8�'�4��(�@���	�ƣ���h]�� ��g�%�|�_�w�}�����ԓ�F9�� 1��U��}�0�
� �a�m�����ƿ�_9��G_�� ��d�%�|�_�w�}�����Փ�F9��1��U��}�8�
�
�"�k�E���Y����@��C�����m�
�g�n�w�}��������U��_��G��u�&�9�!�'�o��������U��[��Gʭ�'�4�
�:�$��ށ�P���F��[1��ߊ� �m�b�%�w�`�_���&˹��lP��h����&�9�!�%��(�O���	����F�D�����
�0�:�2�9�;�(��&���F��T�����m�
�g�:�w�8�(���O�֓�O��N�����!�%�
� �`�h����D�ή�\
��p+�� ���c�
� �`�e�-�W���Y����l��h��B���%�|�_�u�w�8�(���N����Q��G\��H���8�
�
� �a�k�����ƿ�_9��GX�� ��`�%�|�_�w�}�����ޓ�F9��[��G��u�!�%�g��(�F��&����]��R�����3�
�e�l�'�t�}���Y����G��h��D��
�g�i�u�5�2�(��� ����P��Q��C؊�g�:�u�6�'�h��������U��G�U���&�9�!�%�1��O܁�K�����h��Dي�0�:�2�;�1��@؁�KӞ����T�����d�d�n�u�w�.��������D��R1�����
�
�4�!�1��@���	�����h�����0�!�'�'�$�'�_���������Z1�����"�<�0�4�$�:�(ށ�����9��B�\��u�u�&�1��3�(�������R��P ��*���d�d�
�f�k�}�W���Y����lV��1��E��
�
� �d�g��Dϩ�����P��h��D��
�g�e�u�w�l�^ϻ�
��ƹF�N�����;�!�9�f��m�G��I���F��S�����
�'�!�
�$�4��������U��Y�����h�&�1�9�0�>�����ξ�@�������1�&�1�
�9��(�������@��h��D��
�f�y�g�~�W�W���
����]��h�����&�<�;�g�1��@���	���l�N��Uʥ�e�b�
�
�o�k�C���&����l��@��U¼�8�a�3�
�`�j����P���A�R��U���u�u�u�4��2�����ד�V��^����u�&�8�<�#�� �������Z��T��*���d�c�
�d�k�}��������E��X�����0� �&�2�2�u��������l��C�����;�g�3�
�`�d����J���9F������!��"�<�2�<����&����Q��G]��H�ߊu�u�u�u��o�D���I����9��h_�F���u�=�;�}�4�-�(���H����CT�N��R��u�9�0�_�w�}�W���	����@��A]��D��e�e�n�u�w�)���&����A��h��C���%�u�h�}��e����&����CT��EN�����0�e�1�8�%�<�(�������9��UךU���8�d�3�
�e��E��Yۉ��A ��@1��*��
�g�:�u�2���������lU��h�N���u�!�%�
�"�k�O���Y���G��]�����2�;�3�
�`��EϦ�Ӈ��P	��C1��D��n�u�u�!�'����L����[�U�����e�1�8�'�6��F���&����CT��EN����
� �c�c�'�t�}���Y����V��B1�E���u�h�&�1�;�:��������A��M�����;�1�$�
�$�4��������9��B�\��u�u�!�%�f����A����[�Y�����<�
�
� �c�m�����ƭ�l��D��ۊ�|�_�u�u�:��E���&����CT�
N�����d�3�
�l��n��������]��[��D��u�u�!�%�f����O����[�D�����d�'�2�d�a�}����	����@��A_��\�ߊu�u�8�
�c�;�(��&���FǻN��U���
�4�g�d�`�0����&����CU��_��]���0�3�:�
��2�(���N�ד�N��S��D���0�&�u�u�w�}�WϮ�/����@9��h��B���%�n�u�u�w�}����Hƹ��lW��1��U��&�1�9�2�4�+����Q����I��^	��¥��9�
�
�"�d�F���P����]ǑN��U���!�%�d�
�"�l�F܁�H���@��[�����6�:�}�0�>�8�����μ�e��hZ��B���
�g�
�f�{�i�^�ԶY���F��Z��B���
�e�f�%�w�`��������l��C�����/�}�<�;�3�-�!���&����l^��h�Y��|�_�u�u�w�}����H˹��lW�� 1��U��&�1�9�2�4�+����Q����I��^	��¥��9�
�c�1��B؁�J����O��=N��U���u�8�
�l�1��G���	�����h�����0�!�'�'�$�'�_�������]9��O1��#���a�|�_�u�w�)��������9��R��W���"�0�u�!�'�d����OĹ��[��G1�����9�f�`�u�;�8�U���s���F�C��Gڊ� �d�g�
�f�a�W���&����P9��T��]���<�0�&�2�2�u�(���K����A��W�\��|�n�_�u�w�}�W���&�ד�F9��^��D��u�!�
�:�>�����۔��Z��D�����
�
�
�0��d�G��L����9F���*���3�
�d�b�'�}�J���
����U��]�����:�u�%�6�9�)����H��ƹF��Z��F���
�g�b�%�w�`�}���Y���G��[�� ��a�
�f�"�2�}��������U��\�����|�h�r�r�w�1��ԜY���F��G1�*���d�a�
�f�]�}�W���&�ғ�F9��X��G��u�<�;�2�f�;�(��M����K	��V�����
�#�
�|�]�}�W���&�ӓ�F9��1��U��%��9�
��(�F���	����K�
�����e�n�u�u�#�-�Eف�����9��R�����9�
�d�3��i�D���Q����\��XN�\�ߊu�u�8�
�`�;�(��I����[�^�����3�
�a�m�'�}����	����@��A_��\�ߊu�u�8�
�o�;�(��N����[�L�����}�8�
�
�"�h�@���Y�ƭ�l��D��ي�|�0�&�u�g�f�W�������l ��Y�����h�w�w�"�2�}�����Ϊ�C9��d����l��f�3��h�(��Y�ƿ�T�������!�9�f�
�~�}����[����F�C��Fڊ� �d�d�%�w�`��������U��[��G��u�:�;�:�f�t�}���Y���� R��B1�B���u�h�}�:�;�%�2�������l ��X�����u�:�9�-�����I����S��G\����u�u�u�8��j����&����P��G_��Hʦ�1�9�2�6�!�>����������Y�����g�
� �d�b��D��M����9F���*���3�
�f�
�f�a�W���&����|��]��#���
�e�
�g�f�}�W�������V�=N��U���u�8�
�l�4�.�(���H����CW�
N�����2�6�#�6�8�u����ە��]��Q�����4�0��'�4�(���&����A��W�\��|�n�_�u�w�0�(�������9��R��������!�f�h�!���&����CT�N�����u�f�n�u�w�)��������9��R��W���"�0�u�!�'�d����OĹ��[��G1�����9�f�c�u�;�8�U���s���G��_�� ��a�%�u�h�1�-�9���6���� S��h��A���%�}�l�1� �)�W��B�����hZ�����g�d�%�u�j�-�!���&�֓�F9��]��G��u�:�;�:�f�f�W�������9��h_�D���u�h�_�u�w�}�W�������l
��1��3����u�=�;��/����&����l ��\�*��e�u�u�d�~�8����Y���F��Z��A���
�g�d�%�l�}�WϪ�	����U��Z�����h�_�u�u�w�}��������EU��^�E��u�=�;�}�9�8����&����lW�� 1��]���h�r�r�u�;�8�}���Y���G��Z�� ��f�
�a�_�w�}����&����W��N�U���
�:�<�
�2�)�Ǭ�
����F��P ��]���4�&�2�
��(�E���	���O�=N��U���
�f�3�
�g�j����D�ή�\
��p+�� ���c�
� �`�e�-�W�������t#��B��Cڊ� �`�b�%�~�W�W�������l ��[�*��i�u�-�
�#���������F��W��*Ҋ� �d�c�
�d�n�W���Y����G	�UךU���8�
�`�3��k�C���Y����K��C1�����!� �!�'��o�!�������
Q��F�U���u�:�;�:�g�f�W�������9��h_�@���u�h�3�%�4�����*����G��h[��#���3�
�c�m�'�u�F��Hӂ��]��G�U���!�%�`�
�"�l�Dց�M���U��T������'�6� �2�i�(���&����P��G]��Dʱ�"�!�u�m�l�}�WϪ�	����U��[�����h�3�%�6��<��������A��1��M���
�`�b�%��l��������]ǻN�����l�3�
�c�d�-�W������G9��D�����!�'�
�g��e����L�ѓ� N��
�����g�|�_�u�w�0�(�������
_��N�U���
�!��&��)��������l0��h��D��
�f�f�u�8�3���P���F��G1�*���d�g�
�a�k�}��������V9��E�� ���`�
�
�
�"�l�Eׁ�J����W	��C��M��u�u�!�%�a����M����Z�Q�����4�0��'�4�(���&����U��\�����d�1�"�!�w�l�L���YӒ��lP��B1�L���u�h�}�0�$�:��������9����U���6�;�!�9�f�l�L���YӒ��lQ��B1�Lފ�a�i�u�
�6�o�D܁�����
9��]����!�u�g�n�w�}����A����W��G\��H���w�"�0�u�#�-�N���&����CR������!�9�f�b�w�1����[���F��G1�����c�
�a�i�w�u��������F��Z�� ���g�%�u�u�8�1����6����V��B1�B���|�s�7�:���G���&����U��\��G��u�u�!�%�1��C܁�K���W�@��U¦�2�0�}�;�6�-����/���@��R
�����;�!�9�f��t�W�������l�N�����3�
�c�
�e�a�Wǭ�����l��h_�@ʭ�'�4�
�:�$��ށ�P���F��C1��*��
�g�i�u�f�}����Q����T����#���4�
�&�<�9�;�(��&���F��D�����-�
��-�"��Aց�&¹��lU��h�\ʰ�&�u�e�n�w�}��������lW��B1�A���u�h�}�<�9�4�(ށ�����^��Y
�����3�
�b�
�e�f�W�������U
��h_����� �b�d�%�w�`�_���J����_��G\��ʥ�f�
�
� �a�m����s���F��E�����3�
�g�b�'�}�J�������VU��^1��*��d�%�u�;�w�.��������
9��UךU���;�0�3�:����������
9��R��]���0�3�:�
��(�F��&����\��G1�����9�d�d�n�w�}��������lU��B1�A܊�g�i�u�7�:�/����¹��lW��1��U���u�&�0�
��(�F��&���9F������:�
�
�:��(�F��&���F��Y
�����
�
� �d�c��EϦ�Ӈ��P	��C1��D��n�u�u� �3�/����M����R��h�I���7�8�'�0�n�4�(���H����CT��Y
�����
�
� �d�g��D��Y����]��Q��*ފ�:�
� �d�n��E��Yۓ��V��X��*���d�m�
�g�/�/��������_��G�U��� �1�'�9� �;�(��&���F��R	����� �g�l�%�w�3�W�������9��Q��Eފ�g�n�0�1�5�5���