-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ���d���}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e�'�3�4�'�<�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y����C9��T��;ʆ�����]�}�W���&����R
��V1��*���u�u�����0���s���C9��E�����o��u����>���<����N��
�����e�n�u�u�'�l��������C9��SN�<����
���l�}�WϮ�K����Z	��N��U���
���
��	�%���Hӂ��]��G�U���%�g��'�8���������}F��s1��2���_�u�u�
����������\��b:��!�����
����_������\F��d��Uʥ�a��!�8�9��(߁�	����\��b:��!�����n�u�w�-�C�������T9��N�:���������4���Y����W	��C��\�ߊu�u�
�
��4�����ד�C9��SN�:��������W�W���&ƹ��U9��C��U���������4���Y����W	��C��\�ߊu�u�
�
�2���������WF��~ ��!�����n�u�w�-�A�������T9��N�:���������4���Y����W	��C��\�ߊu�u�
�
��4�����֓�C9��SN�:��������W�W���&Ź��G��Y	��*���u� �u����>���<����N��
�����e�n�u�u�'�k�5�������V9��V�����u� �u����>��Y����l^��h:�����0�e�o����3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���&����^��h��*���#�1�o����3���>����F�G1��6���8�;�
�
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���YӖ��l%��^�����d�4�
�9�w�}�"���-����t/��=N��U���`��6�:�w�}�"���-����t/��a+��:���b�1�"�!�w�t�}���Y����l5��C�����9�u�u� �w�	�(���0���9��dװ���<�0�!�'�w�8����Ӌ��u$��t(��Eʼ�u�u�u�4�#�4����:����t#��e/��:�����o����L���YӇ��A��C��:���������9����Ʈ�[��N�����0�!�'�u�$�}�W���A����%��h^�����%�g�d�
�{��$���)����j6��T��=��������	�FÖ�*����f2��~6��H����
�� ���#Ҧ�N����P
��Z��Y���
�� �
���J��I����J��d1��%�����h�!�2�.�?���*����)��
\�@��`�y��
���6��M߮��l5��h:��H���0������:��1����j(��d>��Y���
��
��f�h�[���&����3��X���u�u�6�;�#�3�W�������l
��^��U����
���w�`�P���s���P	��C��U���6�;�!�9�0�>�G��*����|!��T��R��_�u�u�:�$�<�Ͽ�&����GW��D��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����]ǻN�����4�!�4�
��.�E������5��h"��<������}�n�9� ���Y���F�^�E��e�e�e�e�g�m�L���YӅ��@��CN��*���&�f�3�8�e�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�n�u�u�4�3����Y����g9��1����o������!���6���
F��@ ��U���o�u�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'��(���&����F��d:��9�������w�l�W������F��L�E��e�e�e�e�g�m�G���s���P	��C��U����
�!�
�$��W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��e�e�w�_�w�}��������C9��h��*���
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�����u�:�&�4�#�<�(���
�ޓ�@��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I��ƹF��X �����4�
��&�n�;���Cӵ��l*��~-��0����}�l�1� �)�W���C���V��^�E��e�e�e�e�l�}�WϽ�����GF��h=����
�&�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E���_�u�u�:�$�<�Ͽ�&����GW��Q��D���u��
����2���+������Y��E���h�w�e�e�g�m�F��I����V�=N��U���&�4�!�4��	���&����W�=��*����
����u�NϺ�����O�
N��E��e�e�e�e�g�m�G��B�����D��ʴ�
��&�d��.�(��Cӵ��l*��~-��0����}�l�1� �)�W���C���V��^�E��e�e�e�e�l�}�WϽ�����GF��h=����
�&�
�f�m��3���>����v%��eN��Lʱ�"�!�u�|�m�}�G��I����V��^�E��n�u�u�6�9�)����	����@��h��*��o������!���6���
F��@ ��U���o�u�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'��(���O����lW��N��1��������}�F�������V�S��E��d�e�e�e�g�m�G��[���F��Y�����%��
�!�`�;���Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�e�e�u�W�W�������]��G1��*���m�3�8�d�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�E��w�_�u�u�8�.��������l��1����u�u��
���(���-���_��X����u�h�w�d�g�m�G��I����V��UךU���:�&�4�!�6��#���Kù��^9��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I��ƹF��X �����4�
�:�&��+�E��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������!�4�
�:�$��ށ�Y�Ɵ�w9��p'��#����u�e�1� �)�W���C���]ǻN�����4�!�4�
�8�.�(���K���5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��2�����ԓ�\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����W��UךU���:�&�4�!�6�����&����l^�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
���� T��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��h/��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�D���_�u�u�:�$�<�Ͽ�&����G9��\��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�D��w�_�u�u�8�.��������]��[�*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��d�e�w�_�w�}��������C9��Y����
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�d�d�w�]�}�W���
������T�����f�
�e�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�d�e�g�f�W�������R��V�����
�#�
�u�w�	�(���0����p2��F����!�u�|�o�w�m�L���YӅ��@��CN��*���&�
�#�g�f�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�F���s���P	��C��U���6�;�!�9�e�m�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���I��ƹF��X �����4�
�:�&��+�E��Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�c�w�2����I����D��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����]ǻN�����4�!�4�
�8�.�(���M���5��h"��<������}�d�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����W��d��Uʶ�;�!�;�u�'�>��������F��d:��9�������w�k�W������F��L�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lW��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��_�N���u�6�;�!�9�}��������EU��(��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��_�D���_�u�u�:�$�<�Ͽ�&����G9��\��3��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�D��d�n�u�u�4�3����Y����\��h��G��u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��Y����
��o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�d�d�e�l�}�WϽ�����GF��h�����#�g��d�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�F��I����V��d��Uʶ�;�!�;�u�'�>��������F��d:��9�������w�k�W������F��L�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������U��N��1��������}�F�������V�S��E��e�d�e�d�u�W�W�������]��G1�����9�d�
�c�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����W��d��Uʶ�;�!�;�u�'�>��������u#��N��1��������}�F�������V�S��D��d�d�d�e�u�W�W�������]��G1�����9�d�
�`�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��d��Uʶ�;�!�;�u�'�>�����Г�\��c*��:���
�����}�������	[�^�E���_�u�u�:�$�<�Ͽ�&����G9��1�U����
�����#���Q�ƨ�D��^��O���d�e�d�w�]�}�W���
������T�����d�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����]ǻN�����4�!�4�
�8�.�(���K���5��h"��<������}�f�9� ���Y���F�^�E��e�d�n�u�w�>�����ƭ�l��D�����d�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�d�n�w�}��������R��X ��*���d�e�o����0���/����aF�N�����u�|�o�u�g�m�G��I���9F������!�4�
�:�$�����I����g"��x)��*�����}�f�3�*����P���V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g��}���Y����G�������!�9�d�
�g�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��L�U���6�;�!�;�w�-��������9��N�&���������W��Y����G	�N�U��d�d�d�e�g��}���Y����G�������!�9�d�
�a�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��L�U���6�;�!�;�w�-��������9��T��!�����
����_������\F��T��W��e�e�d�e�g�f�W�������R��V�����
�#�g���g�$���5����l0��c!��]��1�"�!�u�~�g�W��H����W��L�U���6�;�!�;�w�-��������9��T��!�����
����_������\F��T��W��e�e�d�e�f�f�W�������R��V�����
�#�g���g�$���5����l0��c!��]��1�"�!�u�~�g�W��H����W��L�U���6�;�!�;�w�-��������9��q(��3�����u�u���8���&����|4�]�����:�e�u�h�u�l�F��H����W��_�D��d�d�d�d�f�l�F��H����W��_�D��u�u�6�;�#�3�W�������l
��1�Oʆ�������8���H�ƨ�D��^��O���e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)����H����g"��x)��*�����}�u�8�3���Y���V��^�W�ߊu�u�:�&�6�)��������_��h]��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�l�L���YӅ��@��CN��*���&�
�#�g���Mύ�=����z%��r-��'���d�1�"�!�w�t�M���H����W��_�N���u�6�;�!�9�}��������EW��V��U���
���
��	�%���Hӂ��]��G��H���e�e�e�d�g�m�L���YӅ��@��CN��*���&�
�#�a���1���Y����)��t1��6���u�g�u�:�9�2�G���D����W��_�D��d�d�d�d�f��}���Y����G�������!�9�g�
�w�}�#���6����e#��x<��G���:�;�:�e�w�`�U��I����V��^�E��e�e�w�_�w�}��������C9��Y����
��u�u���8���&����|4�_�����:�e�u�h�u�l�F��I����]ǻN�����4�!�4�
�8�.�(���K����	F��s1��2������u�f�}�������	[�^�E��e�d�w�_�w�}��������C9��Y����
�b�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�d�d�d�l�}�WϽ�����GF��h�����#�m�f���g�$���5����l0��c!��]��1�"�!�u�~�g�W��H����W��_�D��n�u�u�6�9�)����	����@��A\��B����u�u����>���<����N��
�����e�u�h�w�f�l�F��H����W��_�D���_�u�u�:�$�<�Ͽ�&����G9��Z��E��e�o�����4���:����T��S�����|�o�u�d�g�m�G��I����V��^�E��u�u�6�;�#�3�W�������l
��1��3���o������!���6���F��@ ��U���o�u�e�d�f�l�F��H����D��N�����!�;�u�%�4�3����H˹��V��N��1��������}�F�������V�S��D��e�e�e�e�g�m�G���s���P	��C��U���6�;�!�9�d��D���Cӵ��l*��~-��0����}�a�1� �)�W���C���V��^�E��e�e�e�d�g�m�F��I����D��N�����!�;�u�%�4�3����J����\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lT��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����W��^�N���u�6�;�!�9�}��������E_��T��!�����
����_�������V�S��E��e�e�e�n�w�}��������R��X ��*���
�u�u����>���<����N��S�����|�o�u�d�f�f�W�������R��V�����
�#�
�u�w�	�(���0����p2��F����!�u�|�o�w�l�G��Y����\��V �����:�&�
�#��}�W���&����p9��t:��U��1�"�!�u�~�g�W��H��ƹF��X �����4�
�:�&��+�B��Cӵ��l*��~-��0����}�a�1� �)�W���C���V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�f�f�g�$���5����l0��c!��]���:�;�:�e�w�`�U��[���F��Y�����%�6�;�!�;�n�C��*����|!��h8��!���}�u�:�;�8�m�W��[����l�N�����;�u�%�6�9�)����K����g"��x)��*�����}�u�8�3���Y���W��d��Uʶ�;�!�;�u�'�>�����Փ�\��c*��:���
�����}�������	[�_�N���u�6�;�!�9�}��������EU��V��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��_�E���_�u�u�:�$�<�Ͽ�&����G9��\��C��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�D��e�n�u�u�4�3����Y����\��h��G��u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��Y����
�`�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�d�d�d�l�}�WϽ�����GF��h�����#�g�f�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�d�e�f��}���Y����G�������!�9�f�
�`�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�f�l�F��Y����\��V �����:�&�
�#�f�m�Mύ�=����z%��r-��'���e�1�"�!�w�t�M���I����V��^�E��e�e�w�_�w�}��������C9��Y�����f�o�����4���:����W��X����u�h�w�d�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�g�m�L���YӅ��@��CN��*���&�
�#�g�`��1���Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���W��_�D��d�d�d�d�f�l�F��H����l�N�����;�u�%�6�9�)���&����V��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��N�&���������W������\F��T��W��n�u�u�6�9�)����	����@��A]��E��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[�*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��d�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�d�w�_�w�}��������C9��Y����
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�e�w�]�}�Wϭ�����R��d1����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����D��N�����<� �0�3�:�8��������@��Y	�U���4�!�<� �2�;��������TF����6���&�u�u�<�9�1��������l�N�����u�%�&�2�4�8�(���
�ד�@��T��!�����n�u�w�.����Y����Z��S
��C������]�}�W�������lV��R�����
�;�&�2�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������lV��R�����
�'�2�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�f�W���
����_F��1�����%�4�4�
�;���������g"��x)��N���u�&�2�4�w��(���&����R9��h��*���2�o�����4��Y���9F������%�d�'�3�:�%��������`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�d�'�3�8�/�-����Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�D�����
�
�0�
�6���������@��N��1�����_�u�w�4����	�ד�V ��V�����1�%�0�u�w�	�(���0����A��d��Uʦ�2�4�u�
��8��������TF��d:��9�������w�n�W������]ǻN�����9�%�g��%�2�(�������g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����9�%�g��%�2�(�������]9��PN�&������_�w�}����Ӗ��l6��^�����9�
�'�2�m��3���>���F�UךU���<�;�9�%�b�/��������l��T��!�����
����_������\F��d��Uʦ�2�4�u�
��8�(�������TF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���&�2�4�u����������C9��S1��*���u�u��
���L���Yӕ��]��G1�����7�!�
�%�!�9����Y�Ɵ�w9��p'��O���e�n�u�u�$�:����	����l��h_�U������n�w�}�����Ƹ�C9��1����e�u�u����>���<����N��S�����|�_�u�u�>�3�Ϲ�	����Q��G\��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u��%�>�������9��P1�E���u��
����2���+������Y��E��u�u�&�2�6�}��������B9��h��*���
�u�u����>��Y����Z��[N��*���
�1�
�g�w�}�8���8��ƹF��^	��ʲ�%�3�
�b��o�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��d1��<��� �
�d�
�2��O��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
�0�
�m�`�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����R��^	������
�!�
�$��W���-����t/��=N��U���;�9�4�
�>�����M����q)��r/�����u�<�;�9�#�-�Fہ�����l��N��1��������}�B�������V�=N��U���;�9�!�%�f�����A���5��h"��<������}�f�9� ���Y����F�D�����8�
�
� �b�j����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���0�
�m�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ɗ�l ��Z�����u��
����2���+������Y��E��u�u�&�2�6�}�E�������F��d:��9�������w�l�W������]ǻN�����9���
�����@����	F��s1��2������u�g�9� ���Y����F�D����� ����%�:�D��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����a�3�
�b��n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���
�m�m�o���;���:����g)��[�����:�e�n�u�w�.����Y����l ��^�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�4��������U�=��*����
����u�W������]ǻN�����9�<�;�2�f�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʼ�;�2�d�'�0�n�A���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���3�
�m�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��W�����m�b�o����0���/����aF�
�����e�n�u�u�$�:��������l �� ]�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&���� ^��T��!�����
����_�������V�=N��U���;�9�!�%�f�m����Lƹ��\��c*��:���
�����j��������l�N�����u�8�
�g��8�(��I����g"��x)��*�����}�b�3�*����P���F��P ��U���
�g�
� �`�d����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N����d�'�2�f�n�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h_�� ��b�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������A��W�U����
�����#���Q�ƨ�D��^����u�<�;�9�%�l����Oʹ��\��c*��:���
�����}�������9F������'�d�'�2�d�m�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����
� �m�`�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��[1�����'�2�f�d�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����@��C��L���
�m�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G\�����f�d�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��h��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ����� S��R	��L��o������!���6�����Y��E��u�u�&�2�6�}����&����W��N�&���������W������\F��d��Uʦ�2�4�u�6�'�����@���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�c�
� �n�j����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���'�2�f�f�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������R��1�����0�
�
�d�1��G���	����`2��{!��6�����u�e�3�*����P���F��P ��U���2�g�4�9�8�8�(ށ�H����lU��N�&���������W������\F��d��Uʦ�2�4�u�4�0�l��������9��h��D��
�f�o����0���/����aF�
�����e�n�u�u�$�:��������l��h�����<�
�0�
�n�k�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��Y	��*���
�0�:�
��l����H�ߓ� F��d:��9�������w�m��������l�N�����u�4�2�d�6�1����
�ԓ�9��P1�@���u��
����2���+����W	��C��\�ߊu�u�<�;�;�-�Nف�H����W��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��k�ށ�����^�=��*����
����u�W������]ǻN�����9�%��9�����Oǹ��\��c*��:���
�����n��������l�N�����u�
�4�g�c�/���O����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʴ�
�<�
�&�&��(���&����F��d:��9����_�u�u�>�3�Ͽ�&����Q��W�Oʗ����_�w�}����ӈ��@��U�����f�b�u�u���8���&����|4�N�����u�|�_�u�w�4�������� 9��h_�C���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����K����T9�� Y��U���
���
��	�%���Y����G	�UךU���<�;�9�1�;�)��������F9��X��F��������4���Y����\��XN�N���u�&�2�4�w�8����&����@9��P1�M���u��
����2���+����W	��C��\�ߊu�u�<�;�;�9��������@9��h_�A���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������]��E��F��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1�%���¹��_9��R��*���`�3�
�b�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��V ��D���9�:�0�
���B�������F��d:��9�������w�m��������l�N�����u�
�4�g�f����N����\��c*��:���
�����j��������l�N�����u�
�4�g�f�����@���5��h"��<������}�`�9� ���Y����F�D�����#�'�9�"�f�;�(��O����	F��s1��2������u�g�9� ���Y����F�D�����#�'�9�"�f�/���I����`2��{!��6�����u�e�3�*����P���F��P ��U���0�3�:�
��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʠ�1�'�9�"�f�/���H����`2��{!��6�����u�e�3�*����P���F��P ��U���0�2�d�3��m�E���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����2�d�'�2�c�l�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h8��G��
� �g�d��n�Mύ�=����z%��r-��'���f�1�"�!�w�t�}���Y����R
��h8��G��
�0�
�e�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������D�����
��&�d��.�(���Y����)��tUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�)���@����lR��N�&���������W������\F��d��Uʦ�2�4�u�<�9�4�(���K����CU�=��*����
����u�W������]ǻN�����9�&�2�7�#�/���J����`2��{!��6�����u�e�3�*����P���F��P ��U���4�g�f�
�"�o�@݁�K����g"��x)��*�����}�f�3�*����P���F��P ��U���4�g�f�
�2��G��Cӵ��l*��~-��0����}�f�1� �)�W���s���@��V�����2�7�!�g�1��D���	����`2��{!��6�����u�e�3�*����P���F��P ��U���&�2�7�!�e�/���L����`2��{!��6�����u�e�3�*����P���F��P ��U���'�
� �g�n��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��T�����2�a�`�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӂ��V��h�����
� �g�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[�����'�&�g�'�0�i�A���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������a�
� �g�g��D��*����|!��h8��!���}�f�1�"�#�}�^�ԜY�ƿ�T�������a�
�0�
�g�j�Mύ�=����z%��r-��'���f�1�"�!�w�t�}���Y����R
��G1�����0�
��&�f�����I����g"��x)��N���u�&�2�4�w�-��������S�,��9���n�u�u�&�0�<�W���	����lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�>�0�D������� F��d:��9�������w�m��������l�N�����u�8�
�d�1��B���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�d�'�2�c�j�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��F���
�c�`�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��1����m�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����^��B1�D݊�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����9��P1�L���u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	�֓�F9��_��G��������4���Y����\��XN�N���u�&�2�4�w�8�(���Lù��T9��Y��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)��������U��N�&���������W������\F��d��Uʦ�2�4�u�0��0�Bށ�����T�=��*����
����u�W������]ǻN�����9�&�9�!�'�o����O�ғ�F��d:��9�������w�m��������l�N�����u�0�
�8�b�����H���5��h"��<������}�w�2����I��ƹF��^	��ʴ�
�<�
�&�&��(���K����lW��N��1�����_�u�w�4��������T9��S1�B������]�}�W�������q9��h-�����'�6� �0�f�e����A�ד� F��d:��9�������w�o��������l�N�����u��6�
�6�8�$�������lW��h��*��a�o�����4���:����T��X����n�u�u�&�0�<�W�������9��P1�G���u��
����2���+����W	��C��\�ߊu�u�<�;�;�-�!���&�֓�V��\�Oʆ�������8���J�ƨ�D��^����u�<�;�9�&�4�(ށ����� R�=��*����
����u�W������]ǻN�����9�!�%�d�g�;�(��O����	F��s1��2������u�e�}�������9F������!�%�d�e�%�:�C��Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����d�d�'�2�c�i�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��@؊�0�
�d�l�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��1����`�u�u����>���<����N��S�����|�_�u�u�>�3�Ϯ�+����G9��V�����d�l�o����0���/����aF�
�����e�n�u�u�$�:����&����_��h��*��a�o�����4���:����T��X����n�u�u�&�0�<�W�������9��P1�B���u��
����2���+����W	��C��\�ߊu�u�<�;�;�-�!���&�ԓ�V��Y�Oʆ�������8���J�ƨ�D��^����u�<�;�9�&�4�(݁�����W�=��*����
����u�W������]ǻN�����9�!�%�d�`�;�(��I����	F��s1��2������u�e�}�������9F������!�%�d�b�%�:�C��Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����d�m�'�2�c�d�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��@ӊ�0�
�d�c�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��1����e�u�u����>���<����N��S�����|�_�u�u�>�3�Ϯ�+����G9��E��A��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����
����9��P1�D���u��
����2���+����W	��C��\�ߊu�u�<�;�;�-�!���&����l ��_�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������V��R	��G��o������!���6���F��@ ��U���_�u�u�<�9�1��������V��c1��Dي�&�
�g�o���;���:���F��P ��U���&�2�7�1�d�h�MϜ�6����l�N�����u�
�4�g�b����N˹��\��c*��:���
�����l��������l�N�����u�
�4�g�b�����K���5��h"��<������}�f�9� ���Y����F�D������6�
�4�2���������W��B1�F܊�f�o�����4���:����U��S�����|�_�u�u�>�3�Ϸ�&����R��d�����0�d�d�'�0�i�E���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*���
�&�$���)�C�������	F��s1��2���_�u�u�<�9�1��������W9�� N�7�����_�u�w�4��������l%��R1����� �0�d�m�1��B���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʼ�
�!��&��)��������9��P1�F���u��
����2���+������Y��E��u�u�&�2�6�}�5���&����l5��B�����a�
�4�!�1��A���	����`2��{!��6�����u�b�3�*����P���F��P ��U���6�
�4�0��/��������l��C1����f�u�u����>���<����N��S�����|�_�u�u�>�3�Ͽ�&����P��h=����
�&�
�`�m��3���>����F�D�����%�&�2�7�3�n�N��;����r(��N�����4�u�0�m�1��A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���m�'�2�a�c�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������[�����:�%�d�c�1��A���	����`2��{!��6�����u�d�3�*����P���F��P ��U���9�
�:�
�8�-�F�������S��N��1��������}�FϺ�����O��N�����4�u�%�&�0�>����-����9��Z1�U����
���l�}�Wϭ�����R��^	�����`�u�u����L���Yӕ��]��C��D���3�
�c�`�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�@���2�a�`�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ʃ�Z��Y
�� ��g�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����lR��h��*��o������!���6���F��@ ��U���_�u�u�<�9�1����&����V9��[��*���
�g�l�o���;���:����g)��]����!�u�|�_�w�}����Ӈ��@��T��*���&�d�
�&��e�Mύ�=����z%��N�����4�u�%�&�0�?���L����|)��v �U���&�2�4�u�#�m�C����ד�F��d:��9�������w�n�W������]ǻN�����9�6�
����%�������l��h��*��a�o�����4���:����U��S�����|�_�u�u�>�3�ϼ��֓�R��V
�����u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����I����
9��N�&������_�w�}����ӄ��lV��Z�����u��
����2���+������Y��E��u�u�&�2�6�}����&����l��E��D��������4���Y����\��XN�N���u�&�2�4�w�(�(߁�K�ߓ�VW�=��*����n�u�u�$�:��������T��h��U����
���l�}�Wϭ�����Q��1�Aӊ�d�o�����4���:����U��S�����|�_�u�u�>�3�ϼ��֓�R��F_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�#�m�C����֓�W��D�Oʆ�������8���Hӂ��]��G�U���&�2�4�u�#�m�C����֓�VV�=��*����n�u�u�$�:�����֓�S��h^�����&�d�o����0���/����aF�
�����e�n�u�u�$�:�����֓�S��h^�����u��
���f�W���
����_F��h^��Aߊ�
�
�0�u�w�	�(���0��ƹF��^	��ʹ�
�
�a�
���F��*����|!��h8��!���}�e�1�"�#�}�^�ԜY�ƿ�T����E��`�0�e�$�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����_��hZ�*���
�1�'�&�g�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����_��hZ�*���
�0�u�u���8���B�����Y�����
�a�
�
��9����H����g"��x)��*�����}�u�8�3���B�����Y�����
�a�
�
��8�W���-����t/��=N��U���;�9�9�
��i�(���&����	F��s1��2���_�u�u�<�9�1����&����V9��S_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�#�m�C����ד�F��d:��9�������w�n�W������]ǻN�����9�<�
�<��/�;���&����T9��N�&���������W������\F��d��Uʦ�2�4�u�%�$�:����&����GW��Q��D���u��
���f�W���
����_F��h��*���
�f�u�u���6��Y����Z��[N��*���
�&�$���)�B�������	F��s1��2���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������T9��R��!���g�
�&�
�n�g�$���5����l�N�����u�%�&�2�5�9�C��CӤ��#��d��Uʦ�2�4�u��4�����*����G��h_�*���f�e�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������^��V�� ��f�
�a�o���;���:����g)��]����!�u�|�_�w�}����Ӂ��l ��Y�����u��
����2���+������Y��E��u�u�&�2�6�}��������l��N��1��������}�D�������V�=N��U���;�9�2�%�1��@؁�I����g"��x)��*�����}�d�3�*����P���F��P ��U���
� �a�b�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��V����� �a�f�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����W9��D��*ۊ� �a�c�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����W9��D��*���a�f�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƥ�V��h��A���%�u�u����>���<����N��
�����e�n�u�u�$�:��������C9��Q��Dي�a�o�����4���:����W��S�����|�_�u�u�>�3�Ϫ�	�Г�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(؁�����l��N��1��������}�A�������V�=N��U���;�9�!�%�f����L����	F��s1��2������u�f�}�������9F������!�%�f�
�"�h�@���Y�Ɵ�w9��p'��#����u�`�1� �)�W���s���@��V�����m�3�
�c��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��X�� ���d�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������9��D�����3�
�m�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h8�� ���b�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����T��B1�F���u�u��
���(���-���W��X����n�u�u�&�0�<�W���&�ԓ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w������ד�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�/����H����W��G_��U���
���
��	�%���Jӂ��]��G�U���&�2�4�u�/�����&¹��lP��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�#�-�D؁�����l��N��1��������}�F�������V�=N��U���;�9�!�%�f�e����L¹��\��c*��:���
�����l��������l�N�����u�8�
�m�1��Bځ�J����g"��x)��*�����}�g�3�*����P���F��P ��U���0� �!�b�1��A܁�H����g"��x)��*�����}�f�3�*����P���F��P ��U���
�
�
� �a�j����Y����)��t1��6���u�`�u�:�9�2�G��Y����Z��[N����c�3�
�d��l�Mύ�=����z%��r-��'���g�1�"�!�w�t�}���Y����R
��1�����m�
�g�o���;���:����g)��_����!�u�|�_�w�}����ӷ��}9��t1�����l�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����V��B1�L���u�u��
���(���-���W��X����n�u�u�&�0�<�W���&�ד�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�5����H����W��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�6��(ف�����l��N��1��������}�B�������V�=N��U���;�9�&�
�:��(�������W��G_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�:��A���&����CW�=��*����
����u�DϺ�����O��N�����4�u�8�
�`�;�(��&���5��h"��<������}�d�9� ���Y����F�D�����8�
�d�
�"�j�N���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����a�
� �b�n�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��C��@ڊ� �b�f�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����G��]�� ��l�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Q��V�����m�
�d�o���;���:����g)��]����!�u�|�_�w�}����Ӓ��lS��Q��Bي�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����U��W��F��������4���Y����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��o�(���A�Փ�F��d:��9�������w�h��������l�N�����u�8�
�c�1��F؁�K����g"��x)��*�����}�u�8�3���B�����Y�����d�3�
�g��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�A���
�f�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������P��B1�@���u�u��
���(���-���U��X����n�u�u�&�0�<�W���&����U��_��G��������4���Y����W	��C��\�ߊu�u�<�;�;�-�%�������U��Y��G��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����S��N�&���������W������\F��d��Uʦ�2�4�u�8��j����O����\��c*��:���
�����}�������9F������!�%�a�
�"�j�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�g�
� �o�n����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*��
� �m�`�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������G_�� ��`�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������9��hY�*��o������!���6�����Y��E��u�u�&�2�6�}���A����G9��D�� ��b�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����e9��Q��Aߊ�g�o�����4���:����W��S�����|�_�u�u�>�3�Ϫ�	����U��[��G��������4���Y����W	��C��\�ߊu�u�<�;�;�)���J����
U��GZ��U���
���
��	�%���Iӂ��]��G�U���&�2�4�u�8�l�F���&����CT�=��*����
����u�FϺ�����O��N�����4�u�:�g�f�;�(��&���5��h"��<������}�f�9� ���Y����F�D�����8�
�f�
�"�d�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����d�6�&�
�"�d�D���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����c�
� �l�`�-�W���-����t/��a+��:���`�u�:�;�8�m�L���Yӕ��]��C��Cي� �l�d�%�w�}�#���6����e#��x<��@���:�;�:�e�l�}�Wϭ�����_"��h��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϭ�����l_��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:�j����I�ד�F��d:��9�������w�m��������l�N�����u�8�
�f��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�c�
� �f�o�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��ي� �d�g�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����C	��h_�����3�
�c�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������hX�����e�l�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƞ�]��h8��*���d�a�
�g�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������l0��h��D��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������]��h�����e�f�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӵ��T��V�����
�
� �d�b��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��e��ۊ�9�
�;�&�d�;�(��N����	F��s1��2������u�g�9� ���Y����F�D�����8�
�m�3��m�F���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����d�4�9�/�%�.�E���&����l��N��1��������}�GϺ�����O��N�����4�u�4�2�f�<��������l ��_�*��o������!���6�����Y��E��u�u�&�2�6�}����A����l ��_�*��o������!���6�����Y��E��u�u�&�2�6�}����@����V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����T��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)��������_��N�&���������W������\F��d��Uʦ�2�4�u�'�4�3�N܁�H����V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�6�:�F�������@9��Q��E���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ����� ^��B1�Fߊ�f�o�����4���:����V��X����n�u�u�&�0�<�W���L����U��_�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�-�Nׁ�H����V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����S��G]��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�l�O���&����l��N��1��������}�GϺ�����O��N�����4�u�8�
��(�F��&���5��h"��<������}�e�9� ���Y����F�D�����
�0� �!�a�;�(��A����	F��s1��2������u�b�}�������9F������8�;��d�1��F���	����`2��{!��6�����u�`�w�2����I��ƹF��^	��ʡ�%�g�3�
�e�h����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N�����3�
�g�e�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��*���d�d�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������R��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����
����G9��D�� ��g�
�d�o���;���:����g)��]����!�u�|�_�w�}����Ӓ��l_��B1�A݊�d�o�����4���:����S��S�����|�_�u�u�>�3�Ϫ�	����U��[�����u��
����2���+������Y��E��u�u�&�2�6�}����I����T��h�Oʆ�������8���K�ƨ�D��^����u�<�;�9�#�-�Fށ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��o����K�ԓ�F��d:��9�������w�n�W������]ǻN�����9�!�%�m�1��E���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�a�3�
�e�j����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N��G���
�g�d�%�w�}�#���6����e#��x<��G���:�;�:�e�l�}�Wϭ�����G��[�� ��l�
�g�o���;���:����g)��_����!�u�|�_�w�}����Ӓ��lW��T��*���d�e�
�d�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������^��1��*��e�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������
9��h_�@���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Mʹ��lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������^��N�&���������W��Y����G	�UךU���<�;�9�!�'�h�(���H����CT�=��*����
����u�DϺ�����O��N�����4�u�
�0�"�)����&����l��N��1��������}�B�������V�=N��U���;�9�!�%�f����Kù��\��c*��:���
�����}�������9F������!�%�d�
�"�l�Cف�K����g"��x)��*�����}�u�8�3���B�����Y�����9�
�
� �f�e�(��Cӵ��l*��~-��0����}�f�1� �)�W���s���@��V�����b�3�
�f�a�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h��D���
�g�o����0���/����aF�
�����e�n�u�u�$�:����&����U��Y�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�,�(���H����CU�=��*����
����u�W������]ǻN�����9�$�
�&�>�3�F���&����l��N��1��������}�GϺ�����O��N�����4�u�8�
�f�;�(��K����	F��s1��2������u�e�}�������9F������%��9�
��(�F��&���5��h"��<������}�d�9� ���Y����F�D�����8�
�
� �f�o�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�
� �d�g��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����
� �d�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���d�`�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G[�� ��d�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����G��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4����
����^��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CW��Q��A���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����V��B1�Gߊ�f�o�����4���:����T��S�����|�_�u�u�>�3�ϭ�����R��B1�@ي�g�o�����4���:����V��X����n�u�u�&�0�<�W���&¹��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����L����R��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��A���&����l��N��1��������}�E�������V�=N��U���;�9�&�9�#�-�D���&����l��N��1��������}�E�������V�=N��U���;�9�!�%�`����@����\��c*��:���
�����}�������9F������!�%�1�8�%�<�(���H����CT�=��*����
����u�W������]ǻN�����9�!�%�3��i�O���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����3�
�a�e�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��D\�� ��l�
�g�o���;���:����g)��_����!�u�|�_�w�}����Ӓ��lW��h��D��
�f�o����0���/����aF�
�����e�n�u�u�$�:�����ד�R��Q��A���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l ��[�*��o������!���6��� F��@ ��U���_�u�u�<�9�1����KĹ��lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�����L�Г�F��d:��9�������w�m��������l�N�����u�0�
� �f�n�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��ۊ� �d�`�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��_�����`�g�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lT��Q��@���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϭ�¹��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'�.�(�������S��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�#�-�D߁�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�4�0�o�!�������
T��N�&���������W��Y����G	�UךU���<�;�9�'��;�(��A����	F��s1��2������u�b�}�������9F������:�
�:�1�f�4����L�ԓ�F��d:��9�������w�m��������l�N�����u�4�2�g�6�1����&����V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9��9�8�(���&����lW��h��D��
�f�o����0���/����aF�
�����e�n�u�u�$�:��������l��h�����3�
�`�c�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h]�����c�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӵ��T��V�����&�3�
�c�a�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��V ��D���9�/�'�&�f�;�(��M����	F��s1��2������u�g�9� ���Y����F�D�����8�
�e�;�#�;�(��O����	F��s1��2������u�g�9� ���Y����F�D�����8�
�g�3��k�O���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�d�
� �f�j�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�b�3�
�a�e����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������l�
�
� �f�l�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
�9�
�;�$�;�(��M����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�d��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʥ�l�
�
� �f�k�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��LҊ�
� �d�a��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�b�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������E��*��� �d�m�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����a��R_�����;�&�g�<�1��A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���2�d�4�9�-�/��������Q��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����U�� \�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)�݁�����9��T��!�����
����_�������V�=N��U���;�9�6�'�.�l��������Q��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�6�:�E�������@9��Y�����
�b�g�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��[�� ��c�
�f�o���;���:����g)��^�����:�e�n�u�w�.����Y����A��1�����b�m�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӵ��T��V�����
�
� �
��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʥ�l�
�
� �f�k�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��F���
�b�m�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����C9��[\��*���d�l�
�f�m��3���>����v%��eN��Bʱ�"�!�u�|�]�}�W�������^��^�� ��e�
�d�o���;���:����g)��^�����:�e�n�u�w�.����Y����ZW��B1�Dي�g�o�����4���:����V��X����n�u�u�&�0�<�W�������]9��Q��M���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����U��\�����u��
����2���+������Y��E��u�u�&�2�6�}�(���K�Г�F9��Y��G��������4���Y����W	��C��\�ߊu�u�<�;�;�)���@����^��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����R��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)��������U��N�&���������W������\F��d��Uʦ�2�4�u�0��0�D܁�����
9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�F���&����l��N��1��������}�F�������V�=N��U���;�9�&�9�#�-�C���&����l��N��1��������}�F�������V�=N��U���;�9�!�%�f�l����A�Փ� F��d:��9�������w�m��������l�N�����u�8�g�b�3�0����&����Q��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'����A����\��c*��:���
�����}�������9F������6�'�,�d�>����Aʹ��\��c*��:���
�����}�������9F������&�9�!�%�a�3����&����l��N��1��������}�GϺ�����O��N�����4�u�8�m�1��N���	����`2��{!��6�����u�e�3�*����P���F��P ��U���'�
�
�:��l����@�֓�F��d:��9�������w�m��������l�N�����u�4�2�g�6�1����&¹��G9��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������V_��^_�� ��f�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����VW��[�����g�8�-�<��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʇ�;�0�
�9��3����¹��l ��W�*��o������!���6�����Y��E��u�u�&�2�6�}��������V��h��D��
�f�o����0���/����aF�
�����e�n�u�u�$�:��������CR��Q��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϰ�����Q��1��*��`�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������U��Y�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	�ԓ�F9��\��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������R��N�&���������W������\F��d��Uʦ�2�4�u�0��0�Cށ�����9��T��!�����
����_�������V�=N��U���;�9�1�9�#�9����
�ד�F9��]��F��������4���Y����\��XN�N���u�&�2�4�w�8����&����@9��Y�����l�a�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӂ��V��h�����
�:�
�d�1��G���	����`2��{!��6�����u�e�3�*����P���F��P ��U���0�2�
�d�1��G���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�g�3�
�g�l����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��
�����
�;�&�e�>����Oƹ��\��c*��:���
�����}�������9F������7�8�'�0�`�9��������l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}��������]9��Q��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϼ�����
Q��1��*��m�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����R��P ��*���
� �g�a��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G_�����e�c�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��^�� ��c�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}��������U��V�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����S��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)��������^��N�&���������W������\F��d��Uʦ�2�4�u�0�2�8�(�������G9��h\�@���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������V��h^�����
� �g�e��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��Z�����3�
�d�`�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h]�����d�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӂ��V��h�����<�3�
�e�o�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E����
�0�:�2�9�4����H�ד�F��d:��9�������w�m��������l�N�����u�<�;�4�$�:�(���K����CU�=��*����
����u�W������]ǻN�����9�7�8�'�2�j����&����l��N��1��������}�GϺ�����O��N�����4�u�;�0�1�2�(���K����CT�=��*����
����u�W������]ǻN�����9�:�0�3�8����Hƹ��\��c*��:���
�����}�������9F������&�2�
�&�>�3��������R��N�&���������W������\F��d��Uʦ�2�4�u�8�c�;�(��I����	F��s1��2������u�g�9� ���Y����F�D�����'�0�2�
�����J˹��\��c*��:���
�����}�������9F������!�%�f�
�"�o�@ف�K����g"��x)��*�����}�u�8�3���B�����Y�����9�
�
� �e�k�(��Cӵ��l*��~-��0����}�f�1� �)�W���s���@��V�����8�c�
�0�8�:����&����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�o�(���K����CU�=��*����
����u�DϺ�����O��N�����4�u�'�0�0����LŹ��\��c*��:���
�����}�������9F������&�9�!�%�b�;�(��@����	F��s1��2������u�g�9� ���Y����F�D�����8�`�3�
�e�i����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���g�
� �g�f��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��G1��؊�
� �
� �e�k�(��Cӵ��l*��~-��0����}�f�1� �)�W���s���@��V�����8�g�
� �e�d�(��Cӵ��l*��~-��0����}�f�1� �)�W���s���@��V�����2�
�
�d�1��E���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�d�3�
�e�l����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������&�3�
�g�c�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��D�����f�
�0�:�0�3����K�ԓ�F��d:��9�������w�m��������l�N�����u�0�
�8�c����Mƹ��\��c*��:���
�����j��������l�N�����u�0�
�8�c����O����\��c*��:���
�����}�������9F������!�%�d�3��o�O���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�a�
� �e�j�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��#���
�e�8�-�1��E���	����`2��{!��6�����u�d�w�2����I��ƹF��^	��ʦ�9�!�%�a�1��E���	����`2��{!��6�����u�d�w�2����I��ƹF��^	��ʳ�%�!�'�g�e�i�!���&����l��N��1��������}�F�������V�=N��U���;�9�%��;��@���&����l��N��1��������}�F�������V�=N��U���;�9�%��;��@���&����l��N��1��������}�D�������V�=N��U���;�9�!�%�f�o����J�֓�F��d:��9�������w�e��������l�N�����u�8�
�a��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʧ�g�3�
�f�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h��G���
�f�c�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������Q��Q��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϯ�&����T��h��G��
�g�o����0���/����aF�
�����e�n�u�u�$�:����&����lT��Q��F���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l ��]�*��o������!���6��� F��@ ��U���_�u�u�<�9�1����H�Փ�F9��^��F��������4���Y����\��XN�N���u�&�2�4�w�0�(�������P��N�&���������W������\F��d��Uʦ�2�4�u�
�2�(���&����U��W�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�3��������F9��Z��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������W��N�&���������W������\F��d��Uʦ�2�4�u�-������&����_��h8�� ���b�&�3�
�c�k����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N�����<�3�
�a�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E�����g�3�
�a�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��B���
�a�m�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������lU��^1��*��f�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������T��h
�����;�<�3�
�c�n����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����G���1�8�'�4��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʠ�1�'�9�"�e�;�(��J����	F��s1��2������u�g�9� ���Y����F�D�����#�'�9�"�e�;�(��N����	F��s1��2������u�g�9� ���Y����F�D�����8�d�
� �e�e�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����0�<�<�
�"�o�@ׁ�K����g"��x)��*�����}�u�8�3���B�����Y�� ���'�9�"�g�9�)����M�ߓ�F��d:��9�������w�m��������l�N�����u�
�4�g�e���������9��T��!�����
����_������\F��d��Uʦ�2�4�u�
�6�o�F���&����l��N��1��������}�E�������V�=N��U���;�9�!�%�f�k����L�ѓ� F��d:��9�������w�m��������l�N�����u�8�
�m�1��B���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
��-� ��?��������F��1�����`�b�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�C9��d�����&�9�!�
�6�(�(���H����R��h�Oʆ�������8���K�ƨ�D��^����u�<�;�9�1�-�6���6����Q��B��#���0�l�
�
�"�o�C܁�J����g"��x)��*�����}�f�3�*����P���F��P ��U���
� �g�`��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��X��2��� �
�'�4�2���������l ��[�*��o������!���6�����Y��E��u�u�&�2�6�}��������F��E�����'�� �9�f�;�(��L����	F��s1��2������u�g�9� ���Y����F�D�����:�9�-���)�0�������A9��B�����
�a�c�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��Y�� ��b�
�f�o���;���:����g)��_�����:�e�n�u�w�.����Y����_��B1�Cي�a�o�����4���:����T��X����n�u�u�&�0�<�W���N����S��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����W��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�<�:�n�(���&����T��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�e�(���K����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�d����O�ӓ�F��d:��9�������w�m��������l�N�����u�0�
�8�f�l��������U��\�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	����W��E	��*���g�a�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƪ�C9��S�����`�e��3��k�N���Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����;�1�
�0�:�h�A�������^��N�&���������W��Y����G	�UךU���<�;�9�3�'�3��������W��h��G��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������]��B1�MҊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���*����F9��]��F��������4���Y����W	��C��\�ߊu�u�<�;�;�2�(���¹��lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�8�����&����W��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�;� �8�F���&����l��N��1��������}�E�������V�=N��U���;�9�3�%�9�9�(�������l0��B1�C؊�g�o�����4���:����T��S�����|�_�u�u�>�3�ϰ�����l ��Y�*��o������!���6���F��@ ��U���_�u�u�<�9�1�����ӓ�F9��_��F��������4���Y����W	��C��\�ߊu�u�<�;�;�3� ���M����Q��h�Oʆ�������8���K�ƨ�D��^����u�<�;�9�9�*��������S��N�&���������W��Y����G	�UךU���<�;�9�;� �8�D�������U�� Y�����u��
����2���+������Y��E��u�u�&�2�6�}����Ź��lT��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�8�$���&����Q��G]��U���
���
��	�%���Mӂ��]��G�U���&�2�4�u�2����&����_��G]��U���
���
��	�%���Y����G	�UךU���<�;�9�%�$�;�(��N����	F��s1��2������u�e�9� ���Y����F�D�����0�
�8�`��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʦ�9�!�%�a�1��O���	����`2��{!��6�����u�g�3�*����P���F��P ��U���4�g�m�3��j�G���Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����9�
�
� �e�h�(��Cӵ��l*��~-��0����}�a�1� �)�W���s���@��V�����a�3�
�m�n�-�W���-����t/��a+��:���g�u�:�;�8�m�L���Yӕ��]��C��Mߊ� �g�f�
�f�g�$���5����l0��c!��]���1�"�!�u�~�W�W���������V��@��
� �g�a��n�Mύ�=����z%��r-��'���a�1�"�!�w�t�}���Y����R
��h8��G��
� �g�d��n�Mύ�=����z%��r-��'���a�1�"�!�w�t�}���Y����R
��Z��C���
�m�f�%�w�}�#���6����e#��x<��G���:�;�:�e�l�}�Wϭ�����G��Y�� ��a�
�d�o���;���:����g)��\����!�u�|�_�w�}����Ӕ��lR��B1�F݊�g�o�����4���:����T��S�����|�_�u�u�>�3�ϸ�	����2��B�� ���%�,�d�a��;�(��M����	F��s1��2������u�d�}�������9F������!�%�m�
�"�o�Aށ�H����g"��x)��*�����}�c�3�*����P���F��P ��U���
���,�"�����	����R��h��G��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������l ��V�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������J)��h#�����,�d�b��1��O���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�%�-� ���)�:�������T��a1��*��a�%�u�u���8���&����|4�[�����:�e�n�u�w�.����Y����K+��c�����9�<�9�
�e��(���K����CT�=��*����
����u�AϺ�����O��N�����4�u�-�
������&����Z��h_�*��� �g�b�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��F��
�g�o����0���/����aF�
�����e�n�u�u�$�:����&����l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}����
����9��h]�M���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����@¹��lU��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�����L¹��lU�� 1��U����
�����#���Q����\��XN�N���u�&�2�4�w�8��������l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}����K���� V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�6�/�(ށ�����9��T��!�����
����_�������V�=N��U���;�9��;�2���������l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}����H����l��X��*���f�m�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�f�3�
�g�l����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���3�
�e�a�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������1��*���f�l�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƨ�_��S1�����f�3�
�e�a�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h ��*���3�
�d�l�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������R��*���3�
�d�`�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������hW�����d�d�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӂ��V��h�����3�
�d�`�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������1��*���f�d�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ʈ�^��RZ�����'�4�
�d�1��F���	����`2��{!��6�����u�e�3�*����P���F��P ��U���g�c�1�8�%�<�(���J����CT�=��*����
����u�W������]ǻN�����9�!�%�f�1��F���	����`2��{!��6�����u�e�3�*����P���F��P ��U���0�3�:�
��(�D��&���5��h"��<������}�w�2����I��ƹF��^	��ʺ�0�3�:�
��(�D��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�a�3�
�f�l����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������
�
�f�3��l�B���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����3�:�
�
�8����NĹ��\��c*��:���
�����}�������9F������%��9�
�g��������� 9��T��!�����
����_������\F��d��Uʦ�2�4�u�
�6�o�E��&����_��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�����IĹ��\��c*��:���
�����}�������9F������'�<�<�
�"�n�F݁�K����g"��x)��*�����}�u�8�3���B�����Y�����&�<�;�l�1��E���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�`�3�
�e�o����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��#���
�f�3�
�e�k����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����;�<�
�
�"�n�Dށ�J����g"��x)��*�����}�u�8�3���B�����Y�����l�
� �f�d��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��T�����3�
�g�`�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W�������4��P�����:�0�
�
�"�n�Bځ�K����g"��x)��*�����}�u�8�3���B�����Y��'���0�
�9�
�2�2�(ځ�����9��T��!�����
����_�������V�=N��U���;�9��;�2���������l ��\�*��o������!���6�����Y��E��u�u�&�2�6�}����N���� T��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��l�݁�����9��T��!�����
����_�������V�=N��U���;�9�1�9�#�9����
�ғ�F9��[��F��������4���Y����\��XN�N���u�&�2�4�w�����K���� T��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�%�8����M���� U��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��O���&����l��N��1��������}�GϺ�����O��N�����4�u�0�0�2�����J���� T��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��e�݁�����9��T��!�����
����_�������V�=N��U���;�9�7�8�%�8�G�������]9��h��F��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������l��X�����
�f�b�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��h��F��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������_	��1��*��l�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������_	��1��*��`�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������l ��]�*��o������!���6�����Y��E��u�u�&�2�6�}��������ZR��B1�Aފ�g�o�����4���:����V��X����n�u�u�&�0�<�W�������D9��Y�����f�c�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӗ��R
��^�����3�
�f�g�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��a��*ي�d�3�
�f�g�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��C��B���
�f�c�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����Z*��X
�����
�f�
� �d�d�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����l�3�
�f�b�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��^"�����&�
�!� �#�/�(��&ǹ��lU��1��U����
�����#���Q����\��XN�N���u�&�2�4�w���������G��C��*��
�
� �f�g��E��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*��
� �f�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�D���
�a�a�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���f�f�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G\�*���:�2�;�3��i�F���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����e�
� �f�e��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����m�3�
�a�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����c�1�8�'�6����Oʹ��\��c*��:���
�����}�������9F������!�%�d�f�1��C���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�c�
�"�n�@ځ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�d�3��i�F���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�`�
� �d�k�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�b�3�
�c�h����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������4�0��'�4�(���L�ғ�F9��Z��G��������4���Y����W	��C��\�ߊu�u�<�;�;�2�(�������lU��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�9�*��������Q��N�&���������W��Y����G	�UךU���<�;�9�;� �8�O���&����l��N��1��������}�D�������V�=N��U���;�9�:�
�8�9�(���J����CT�=��*����
����u�W������]ǻN�����9�:�
�:�3����Jù��\��c*��:���
�����}�������9F������;�"�0�d��(�D��&���5��h"��<������}�f�9� ���Y����F�D�����0��9�e�1��B���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʻ�"�0�d�
�"�n�Cہ�J����g"��x)��*�����}�d�3�*����P���F��P ��U����9�f�3��h�E���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����0�d�
� �d�k�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����9�a�3�
�b�m����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����d�
� �f�o��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�� ��&���m�3�
�`�o�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��Y����
� �f�l��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��Z��Cފ� �f�a�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��X�����c�f�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lW��h��F��
�d�o����0���/����aF�N�����u�|�_�u�w�4����	����_��X�����&�3�
�c�f�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��C��D���3�
�c�a�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��*���f�l�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƽ�Z*��C1�����:�
�4�!�1��A���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�g��'�:����������\��h��F��
�f�o����0���/����aF�N�����u�|�_�u�w�4����
����^��Q��B���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ����� 9��h]�L���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������U��W�����u��
����2���+������Y��E��u�u�&�2�6�}��������Q��N�&���������W������\F��d��Uʦ�2�4�u�0��0�A���&����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�i����N�ғ� F��d:��9�������w�n�W������]ǻN�����9�<�
�0�:���������]��X�����3�
�b�c�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��7���!�g�l�3��j�C���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�������g��#�o�E���&����l��N��1��������}�D�������V�=N��U���;�9�2�%�1��@ށ�����g"��x)��N���u�&�2�4�w�-��������`2��C\�����u�u��
���L���Yӕ��]��V�����1�
�d�b�m��8���7���F��P ��U���&�2�6�0��	��������\��c*��:���n�u�u�&�0�<�W���
����W��]�Oʗ����_�w�}����Ӈ��@��T��*���&�a�3�8�d�g�$���5����l�N�����u�%�&�2�5�9�E��Y�Ǝ�|*��yUךU���<�;�9�4��4�(�������@��Q��A�������W�W���������D�����g�`�u�u���6��Y����Z��[N��*���
�&�$���)�(���&����`2��{!��6�ߊu�u�<�;�;�<�(���&����W��T��:����n�u�u�$�:��������lR��h��Oʆ�����]�}�W�������C9��h��U����
�����#���Q����\��XN�N���u�&�2�4�w�-��������F��u!��0���_�u�u�<�9�1��������W9��T��:����n�u�u�$�:����	����l��hY�Oʗ����_�w�}����Ӈ��@��U
��M���u����l�W�W�������V��ZV��7����
�
�1�!�n����K����9��~=ךU���0�0�<�u�]�}�W���Y���/��r)��N���u�u�u����6���Cӯ��v!��d��U���u�1�;�
��	�W���7����a]ǻN��U���<�d����g�>���>����F�N�����
���u�w��2���Y��ƹF��X��]���u�u�u�6�<�g�>���-����t/��=N��U���u�0�0�u�w��$���5����l�N��Uʱ�;�u�u����;���:����g)��]����!�u�|�_�w�}�W������/��d:��9�������w�n�W������]ǻN��U���0�o��u���8���B���F�
����������4���:����U��S�����|�|�_�u�w�3�W���	����G]Ǒ=N��U���%�;�;�u�o��Fޝ��֓�C��h]����
�u��u�w�:������ƹF�N��1������]�}�W���Y����`2��rN�<�����_�u�w�}�W���I����g.�'��0���n�u�u�u�w�9����0����	F��c+��'���_�u�u�:�#�u�W���Y����Z��N��U���
���
��	�%���Hӂ��]��G�U���u�u�1� �w�}�"���-����t/��a+��:���c�u�:�;�8�m�W��Y����]��X�����n�_�u�u�4�0����Ӌ��u$��t(��E���3�e�d�a�w��W�������Z�=N��U���u�4�4�<�#�}�W���<����9F�N��U���'�&��;�2�g�>���>����F�N��4���0�&�<�!�w�}�9���<���9F������u�u�u�u�4�6�Mϗ�Y����)��tUךU���u�u�0�0�w�}�9ύ�=����z%��N��U���4�1�0�&�w�}�9ύ�=����z%��r-��'���u�:�;�:�g�f�W���Y����VV�'��&������_�w�}�W���I����f2��c*��:���
�����l��������l�N��Uʴ�1�0�&�u�w��$���5����l0��c!��]���:�;�:�e�l�}�W���YӅ��\��yN��1�����_�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u�3�}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY���F��T�� ����
�����#���Q����\��XN�U��u�u�0�1�4�0������ƓF�T�����!�8���f��(߁��֓�S��h^��&���u�2�;�'�4�u�W���Y����R��^
��U������n�w�}�W���8����@��Y	��Oʜ����_�w�}�W�������@1��C��U�����u�n�w�}����Y���F�N�����u��
���L���Y�����R��U��������W�W���Y�ƭ�W��D^��U���������4���Y����\��XN�N���u�u�u�6�g�g�>���-����t/��=N��U���u�e�o����3���>����v%��eN��Eʱ�"�!�u�|�]�}�W���Y����V��T��;ʆ�������8���Hӂ��]��G�U���u�u�6�d�m��W���&����p]ǻN��U���0�u�u����;���:���F�N��U���������!���6���F��@ ��U���_�u�u�u�w�l�Mϑ�-ӵ��l*��~-��0����}�e�1� �)�W���P���F��SN�����0�!�_�_�5�:����Yӄ��lV��Z�� ��6�8�:�0�#�0�1���H����9��Q1��D��_�u�u�0�2�4�W���Y���F�N�����1�=�h�u�e�W�W���Y�ƍ�W��D<�����k�f�_�u�w�}�W�������Z��S�G�ߊu�u�:�!�:�-�_���Y�����S����9�y�u�u�w�}�������R��D�U���u�u�4�1�2�.�W�������lW��1�����&�y�u�u�w�}���D�Ʈ�U9��\�*���y�u�u�u�w�,�W�������lW��1��Y���u�u�u�4�3�8����Gӄ��lV��Z�����0�&�y�u�w�}�WϽ�H���Q��1�Aӊ�0�y�u�u�w�}� ��D�Ʈ�U9��\�*���y�u�u�u�w�9�W�������lW��1��Y���u�u�u�$�w�c����I����
9��UװU���9�
�
�a���(���Y����\��CN��3���d��
�
�#�m�C�����ƹF��R �����4�u�_�u�w�}�W�������[F�]����u�u�u�1�%�.�%������ JǻN��U���1�'�&��3�5�J���P�����CN�����u�u�u�u�4�6�J���	����l�N��Uʧ�&�!�h�u�'�/��ԜY���F��S�����k�9�
�
�c��(߁�����@V�N��U���6�e�h�u�#�m�C����֓�VV�N��U���$�u�k�9���Cځ�&ù��l�N��Uʴ�1�0�&�u�i�1�(߁�Mƹ��9��S�����u�u�u�u�4�l�J����֓�S��h^�����u�u�u�u� �l�J����֓�S��h^�����u�u�u�u�3�}�Iϲ�&ù��9��1��Y���u�u�u�$�w�c����&����V9��F_����u�9�
�
�c��(ށ�Y�Ư�^��R ��ғ��d��
��(�(߁�K��ƹF��R �����4�u�_�u�w�}�W�������[F�]����u�u�u�1�%�.�%������ JǻN��U���1�'�&��3�5�J���P�����CN�����u�u�u�u�4�6�J���	����l�N��Uʧ�&�!�h�u�'�/��ԜY���F��S�����k�9�
�
�c��(ށ�����@V�N��U���6�e�h�u�#�m�C����ד�VV�N��U���$�u�k�9���Cځ�&¹��l�N��Uʴ�1�0�&�u�i�1�(߁�Mƹ��9��S�����u�u�u�u�4�l�J����֓�S��h_�����u�u�u�u� �l�J����֓�S��h_�����u�u�u�u�3�}�Iϲ�&ù��9��1��Y���u�u�u�$�w�c����&����V9��F_����u�3�e�3�>��E���J���� T��h;�Oʶ�8�:�0�!�:��5���?����U��h]����;�
�g�b�w�}��������R�=N��U���u��h�u�{�}�W���YӨ��l5��p+��K��_�u�u�u�w�4�G���=���F��d��U���u�1�;�
��	�W���J��ƹF�N��������h�w�o�}���Y������FךU���u�u�9�u�i�<�(���U���F������k�4�
�&�{�}�W���Yӂ��F�	��*���a�d�%�y�w�}�W�������X��E�� ��d�%�y�u�w�}�WϽ�Y����A��B1�D���y�u�u�u�w�9����GӁ��l ��Y�����_�u�u�3�g�;����K������\��*��o�6�8�:�2�)�ט�;�׏�U9��Q
��*���&�f�;�
�e�j�W�������Z��V�����u�u�u��j�}�[���Y���(��h=��2���k�b�_�u�w�}�W���I����g.�	N�Y���u�u�u�1�9��>���Y���JǻN��U���:�!����`�W��s���C	����U�ߊu�u�u�u�;�}�IϿ�&����9F�N��U���0�u�k�4��.�[���Y�����N��U���
� �a�b�'�q�W���Y����Z��
P����� �a�b�%�{�}�W���YӅ��X��E�� ��b�6�y�u�w�}�WϺ������h��A���%�|�_�u�w�;�G���������Z��*��o�6�8�:�2�)�ט�;�׏�U9��Q����;�
�a�d�w�}��������R�=N��U���u��h�u�{�}�W���YӨ��l5��p+��K��_�u�u�u�w�4�G���=���F��d��U���u�1� �
��	�W���O��ƹF��X�����}�u�u�u�w�9����Gӂ��@��Y1��*��
�e�_�u�w�}�W������W9��D��*���a�f�%�|�]�}�Wϸ�I����K�� ��Cފ�
�f�o�6�:�2����ˠ��W��Q1�����!�f�;�
�c�l�W�������Z��V�����u�u�u��j�}�[���Y���(��h=��2���k�d�_�u�w�}�W���I����g.�	N�Y���u�u�u�1�"��>���Y���OǻN�����8�%�}�u�w�}�WϺ������D�����3�
�m�
�g�W�W���Y�ƨ�F�	N�����2�
�
� �c�k����s��Ɠ9F�C����6�'�0�!�$�<����	����U�������&�4�0�8�4�4����T�����t=�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W�������F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�]�}�W���Y���F�N������3�8�i�w�-�9���
��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m��������l��A�����u�&�<�;�'�2����Y��ƹF��h^�����9�=�
�%�!�9����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1�����4�%�4�4��1�(������R��X ��*���<�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U���}�4�
�:�$�����&���R��^	������
�!�e�1�0�F���Y����l�N��U���u�u�u�u�w�}�WϮ�I����l��_�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����`�|�!�0�w�}�W���Y���F�N��U���u�
�
�0��1����	����l��PN�U���
�0�
�9�?��������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�e�'�1�<����	����R��P �����&�{�x�_�w�}�(߁�����C��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
��8�(�������V�
N��*���&�
�#�g�g�W�W���Y���F��DךU���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�
�
�0��1����	����F��SN�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^���Y����l�N��U���u�u�u�u�w�-�G�������[��E��I���
�
�0�
�;�5�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�d�'�1�0����&����C�������%�:�0�&�w�p�W���	�ד�V ��V�����1�%�0�
�$�4��������C��R�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���A�C�����u�u�u�u�w�;�_������A��N���ߊu�u�u�u�w�}�W���&¹��U9��O1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�0�$�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-��������`2��C\�����d�|�u�=�9�W�W���Y���F�N��U���u�%�d�'�1�0����&����C��R�����:�&�
�:�>��L���Y���F�N��U���u�9�<�u�6���������F��R ��U���u�u�u�u�w�}�W���Y����lW��R�����%�#�1�%�2�}�JϮ�H����l��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����A��Z�����u�&�<�;�'�2����Y��ƹF��h_�����4�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ד�V ��V�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�d�'�1�0����&����O��_�����u�u�u�u�w�}�W���Y����A��Z�����u�h�%�d�%�;����s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
��8��������W9��R	�����;�%�:�0�$�}�Z���YӖ��l6��^�����9�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�ԓ�V��S1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�0�$�W�W���Y���F�N��U���%�6�;�!�;�:���DӇ��P������u�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-��������`2��C\�����d�|�u�=�9�W�W���Y���F�N��U���u�%�g��%�2�(�������A��S�����;�!�9�2�4�m�}���Y���F�N��U���0�&�3�}�'�.����������YNךU���u�u�u�u�w�}�W���Y�Ƽ�9��E��*���#�1�%�0�w�`����)����W9��h��N���u�u�u�u�w�}�W���YӃ����=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�K����Z	��G��U���<�;�%�:�2�.�W��Y����lT��R�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(݁�����l��PN�U���6�;�!�9�d��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N������'�:�
�'�+����Y����l�N��U���u�u�u�u�w�-�E�������C��R������'�:�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����'�3�7�!��-����	����R��P �����&�{�x�_�w�}�(ځ�����G��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(ځ�����G��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�0�
�2�<��������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&���G��d��U���u�u�u�u�w�}�W���YӖ��l��h�����
�9�
�'�0�a�W���&����Q��h�����_�u�u�u�w�}�W���Y���V��^�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����A��U��*���2�4�&�2�w�/����W���F�G1�����7�!�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l��h�����0�u�h�4��2�����ԓ�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
��8�(�������E
��G�����_�u�u�u�w�}�W���Y���C9��E�����
�'�2�i�w��(���&����l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�;���&����	��h�����`�u�&�<�9�-����
���9F������:�
�:�%�$�/���@����Z��G��U���'�6�&�u�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H��r�u�=�;�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���A����lW��N�����u�u�u�u�w�}�W���Y����9��h(��*���%�&�'�2�c�d�K���5����u	��{��*��
�0�
�g�d�W�W���Y���F�N�����}�4�
�:�$�����&���R��^	������
�!�c�1�0�F���Y����l�N��U���u�u�u�u�w�4�(���?����\	��D1����l�i�u�%�4�3����K����F�N��U���u�u�0�1�>�f�W���Y���F��Y
�����u�u�u�u�2�9���Y����]��E����_�u�u�x�6�.��������@H�d��Uʥ�:�0�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��|�!�0�_�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��CV�����|�|�!�0�]�}�W���Y���F�q\�����m�e�i�u�e�;�(��&����F�N��U���u�u�����(���&����Z�f;��*���
� �`�l�'�f�W���Y���F�N�����d�4�9�:�2��(�������
R��S�����d�4�9�:�2��(�������U��UךU���u�u�u�u�w�}����H����l��X��*���'�2�f�`�w�`�%���¹��_9��E��G���
� �d�`��n�}���Y���F�N��'���0�
�9�
�9�.�F���&���� _��R��'���0�
�9�
�9�.�F���&����P��G]�U���u�u�u�u�w�}����K����lU��N�U���%�
� �l�f�-�L���Y���F�N��U���%�'�2�f�a�}�JϷ�����lP��h����u�u�u�u�w�}�W�������A��V�U��<�0�
�
��(�A���	������Y��C���_�u�u�u�w�}�W���Y����T9��P1�D���h�<�0�
��(�C���	������Y��C���_�u�u�u�w�}�W���Y����l��E��F���u�h�%�l��l����H�ӓ�]ǻN��U���u�u�u�u�5�l����J����[��U1�����l�
�f�_�w�}�W���Y���F��1����e�u�h�'�f�;�(��&����F�N��U���u�u�&�9�#�-�@�������F���*���g�
� �m�b�-�L���Y���F�N��U���
�8�g�
�2��N��E�ƿ�_9��G\�����m�
�g�_�w�}�W���Y���F��[1�����'�2�f�g�w�`��������l ��_����u�u�u�u�w�}�W�������V��R	��M��i�u�8�
�e����L����9F�N��U���u�u�u�8��o�(���&����Z�C��D���3�
�c�
�f�W�W���Y���F�N����
�0�
�m�`�a�W���&�ғ�F9��1��N���u�u�u�u�w�}�WϪ�	����A��V�U��!�%�f�
�"�k�F���B���F�N��U���u�8�
�f�%�:�D��Y����^��1��*��
�g�_�u�w�}�W���Y���G��Z�����m�m�i�u�:��C���&����CU��N��U���u�u�u�u�#�-�Aށ����� R�
N����
� �l�b�'�f�W���Y���F�N�����
�0�
�m�e�a�W���&����lS��h����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���K�V�����'�6�&�{�z�W�W�������@F��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���^�Ƹ�VǻN��U���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�d����A���G��=N��U���u�u�u�u�w�<��������]��1��Dߊ�0�
�l�a�k�}����H����l	��D1����
� �d�m��o�}���Y���F�N�����'�0�
�0��m�@��Y����A��h��G���
�g�_�u�w�}�W���Y���W��C�����
�0�
�l�n�a�W�������\��h��D��
�f�_�u�w�}�W���Y���W��C�����&�'�2�f�o�}�JϺ�����l��X�� ��d�
�f�_�w�}�W���Y���F��@�����
�0�
�l�g�a�W����ԓ�l ��Z�*��g�u�:�;�8�o�^�ԜY���F�N��Uʺ�0�3�:�
��8�(��O���\��Q��*ۊ� �g�d�
�e�W�W���Y���F�N��#���
�l�'�2�d�d�W��	����9��h��D��
�f�_�u�w�}�W���Y���C9��[\��*���
�l�f�i�w�����M����R��h����u�u�u�u�w�}�W���&�Փ�V��Y�I���8�
�f�3��h�A���B���F�N��U���u�;�0�3�8��(���&����Z�B �����"�d�3�
�g�i���Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u�z�}����Ӗ��P��N����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��Dڊ�&�
�|�|�#�8�}���Y���F�N�����,�'�2�a�b�}�JϽ�����F9��\��G�ߊu�u�u�u�w�}�W�������W9��E��G���2�a�c�u�j�9��������\��h��G��
�g�_�u�w�}�W���Y���]��^	�����
�0�
�e�g�a�W����ԓ�9��h\�G���}�f�1�"�#�}�D��Y���F�N��U���
�4�g�d��8�(��K���C9��[\��C���
�g�`�%�l�}�W���Y���F������f�
�0�
�g�i�K���&����lU��Q��F���%�n�u�u�w�}�W���Y����Z��^�����e�c�i�u��<�E��&����_��G\��Aʱ�"�!�u�a�l�}�W���Y���F���*��
�0�
�e�f�a�W����ԓ�9��h\�@���}�f�1�"�#�}�D��Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u�z�}����Ӗ��P��N����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��Dӊ�&�
�m�|�w�5����Y���F�N��U�������#�/�(��&����A��\�U��9�
�
�a���(��s���F�N��U���9�
�
�a���(�������lR��N�U���e�a�`�0�g�,�L���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�u�u�x�w�.����	����@�CךU���'�6�&�u�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H��r�u�=�;�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�����c�|�u�=�9�}�W���Y���F������,� �
�d��8�(��K���T��Q��B݊�g�_�u�u�w�}�W���Y�ƪ�l��a����d�'�2�f�g�}�JϹ�	����Q��G\�U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K��D��ʥ�:�0�&�u�z�}�WϮ�����N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W��PӒ��]l�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�i����H�����Yd��U���u�u�u�u�w�4�(���:����`��T����d�'�2�a�e�}�JϷ�&����R��d�����0�d�d�3��h�A���B���F�N��U���u��6�
�6�8�$�������lW��h��*��a�i�u��4�����*����G��h_�*���f�b�
�f�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�4�&�0�}����
���l�N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���|�!�0�_�w�}�W���Y���F��h��3����:�
�l��8�(��J���Z*��^1�����:�
�l�
�"�n�Eց�K���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϿ�
����C��R��U���u�u�%�:�2�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�d�|�#�8�}���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���d�3�8�d�~�t����s���F�N��U���<�8�f�'�0�i�@���Dӏ��CU��B1�Mۊ�g�_�u�u�w�}�W���Y�Ƽ�e��hZ�����a�c�u�h�'��݁�H����S��h����u�u�u�u�w�}�W���&����9��P1�L���h�&�9�!�'�e����O�ѓ�]ǻN��U���u�u�u�u�2����&����V��R�����!�%�e�3��k�F���B���F�N��U���u�0�
�8�b�����H���F��[1�����3�
�c�f�'�f�W���Y���F�N�����d�'�2�a�`�}�JϪ�	����U��W����u�u�u�u�w�}�W������� 9��P1�M���h�!�%�m��(�E��&����F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W������]F��X�����x�u�u�%�8�8����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�d�~�)��ԜY���F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�g�3�8�f�t�^Ϫ����F�N��U���u�%��&�;��(���&����Z�Q�������!��;�4����Kǹ��U��X�����c�1�"�!�w�i�L���Y���F�N��U���0� �!�f�%�:�C��Y����K��z;�����
� �!�%�.�l�@�������R��F�U���;�:�`�|�]�}�W���Y���F�G1�����
�
�0�
�e�l�K�������f*��x��8���<�9�
�g�����Nǹ��S��S�����a�n�u�u�w�}�W���Y����l4��B����
�0�
�d�n�a�W���&����g��C1�����9�
�g�
��(�E��&���F��@ ��U���n�u�u�u�w�}�W���YӖ��R
��^�����d�l�i�u�/��:��� ����~��^��*��
�
� �g�a��E��Y����G	�G�U���u�u�u�u�w�}��������l��hZ�C��u�-�
���$��������_��Y��*���g�b�
�g�b�}��������l�N��U���u�u�u�$�>��(���&����Z�Q�������!��;�4����Kǹ��U��X�����d�1�"�!�w�l�L���Y���F�N��U���!�g�'�2�c�e�W������~3��N!��*���!�%�,�d�`�����A�ғ�N��
�����g�|�_�u�w�}�W���Y���@��C��G���2�a�e�u�j�.����	�ԓ�F9��Z��G�ߊu�u�u�u�w�}�W�������G9��E��A��u�h�3�%�/��#�������G��N1�A���3�
�m�a�'�u�AϺ�����P�=N��U���u�u�u�u�w�4����&����T9�� ^��Hʳ�%�-� ���)�:�������T��a1��*��a�%�}�c�3�*����O��ƹF�N��U���u�u�8�
�b�����H���F��G1�E���
�l�c�%�l�}�W���Y���F���*���
�0�
�d�c�a�W���&����g��C1�����9�
�g�
��(�E��&��� F��@ ��U��n�u�u�u�w�}�W���YӒ��lW��h��*��l�i�u�-���;�������_��[��Gފ�
� �g�c��o�E�������T��d��U���u�u�u�u�w�)���M����lR��N�U���
���,�"�����	����R��h��G��
�g�`�u�8�3���P���F�N��U���u�!�%�d�`�/���A�����h_�*���g�m�
�d�]�}�W���Y���F�C��D���'�2�a�l�w�`��������J)��h#�����,�d�b��1��O���	������Y��@���_�u�u�u�w�}�W���Y����S��E��A��u�h�3�%�/��#�������G��N1�B���3�
�m�a�'�u�EϺ�����T�=N��U���u�u�u�u�w�0�(��&����T��R�����-� ���#���������9��Q��M���%�}�a�1� �)�W��B���F�N��U���u��6�
�6�8�$�������lW��h��*��a�i�u��4�����*����G��h_�*���g�g�
�f�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�4�&�0�}����
���l�N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���|�!�0�_�w�}�W���Y���F��a��*���'�2�a�g�w�`��������l ��]�*��_�u�u�u�w�}�W���Y����_T��h\�����a�d�u�h�'��݁�&�֓�F9��W��F�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�Fف�
����O�C�����u�u�u�u�w�}�W���A����lR��N�U���m�3�
�c�o�-�L���Y���F�N��U���6�
�4�0��/��������l��C1����f�}�|�i�w���������G��C��*��
�4�!�3��k�B���Q����F�B,�����&�
�!� �#�/�(��&����l��hZ�L��u�h� �
�$���������F��Z�����
� �f�d��l�F��Y����q9��h-�����'�6� �0�f�e����&����T��\��I����6�
�4�2���������^��V�����c�`�%�}�~�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߊu�u�x�4�$�:�W�������K��N�����0�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��D���!�0�_�u�w�}�W���Y���N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l�� 1����|�4�1�}�/�)��������U��N�����:�&�
�#��t�^Ϫ����F�N��U���u�!�%�d�b�/���L����Z�C��D���3�
�c�`�'�u�^�ԜY�Ƹ�C9��1����`�}�|�i�w�0�(��&����U��G_��\�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�l�JϿ�&���R��Y�����<�
�1�
�g�t�^Ϫ����F�N��U���u�!�%�d�e�/���I�����h>�����<�
�<�}�f�9� ���Y���9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�}�W�������@��C�����
�a�
�4�#�/���J����W	��C��\��u�e�e�e�l�}�WϪ�	����l��hZ�M��u�:�;�:�e�}�J���I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�L�ԜY����� ��ʦ�4�0�}�%�������Ƹ�VF��V�����<�0�u�x�w�}����*����l��^	�����u�u�'�6�$�}����*����F��h��U���&�2�7�1�f�d�W�������l ��X�*��_�u�u�0�>�W�W���Y�Ư�@��G1��*���u�&�u�u�w�}�W�������R��c1��D���8�e�h�u�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN��´�
�<�
�1��m�^�������F�N��U���u�u�u�u�6��$������R��c1��G���8�d�_�u�w�}�W���Y���V
��=N��U���u�u�u�u�w�}�W���7����^F���&���!�
�&�
�l�}�W���Y���F���U���_�u�u�u�w�}�W���Ӈ��`2��C\�����u�k�_�u�w�}�W���Y���R��d1����u�%��
�#�����B���F�N��U���;�4�
��$�n����K���9F�N��U���u�u�u�%������DӇ��`2��CZ�����n�u�u�u�w�}�Wϩ��ƭ�l5��D�����f�h�u�u�w�}�W���Y�����y=�����h�4�
��$�h����M���F�N��Uʢ�0�u�%���)�(���&���l�N��U���u�u�u�4������E�ƭ�l5��D�����`�_�u�u�w�}�W�������C9��h��*���
�u�k�_�w�}�W���Y���F��h �����i�u�%���)�(���&��ƹF�N��U���=�;�4�
��.�@������FǻN��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W�������R��c1��M���8�b�h�u�w�}�W���Y���F��G1��*���u�h�4�
��.�N�������F�N��U���"�0�u�%���ց�
����X�N��U���u�u�u�u�6��$������R��c1��Dڊ�&�
�n�u�w�}�W���Yӑ��]F��h=����
�&�
�u�i�W�W���Y���F�N��*���3�8�i�u�'��(���H����lW��=N��U���u�u�u�=�9�<�(���
����U��^��K�ߊu�u�u�u�w�}�W���	����U��S�����
�!�g�3�:�l�L���Y���F���ʴ�
��&�d��.�(��D��ƹF�N��U���u�u�%���.�W������l��1����n�u�u�u�w�}�Wϩ��ƭ�l5��D�*���
�g�h�u�w�}�W���Y���F��G1��*���u�h�4�
��.�Fہ�
����l�N��U���u�"�0�u�'��(���M����lW��
P��U���u�u�u�u�w�}����*����Z�V��!���d�
�&�
�c�W�W���Y���F��R �����
�!�`�3�:�l�W���s���F�N��U���4�
��3�:�a�W���*����P��D��@�ߊu�u�u�u�w�}��������l��1����u�k�_�u�w�}�W���Y���R��d1����u�%��
�#�j����H��ƹF�N��U���=�;�4�
��.�F؁�
����[�=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Q����P	��h��F��
�g�h�4��2����¹��O�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�l�1�0�F��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�Fׁ�
����l�N��U���u�u�u�0�3�4�L���Y���F���ʴ�
��&�d��.�(��D��ƹF�N��U���u�u�%���.�W������l�� 1����n�u�u�u�w�}�Wϩ��ƭ�l5��D�*���
�m�h�u�w�}�W���Y���F��G1��*���u�h�4�
��.�E߁�
����l�N��U���u�"�0�u�'��(���I����lW��
P��U���u�u�u�u�w�}����*����Z�V��!���d�3�8�e�]�}�W���Y���D�������h�u�_�u�w�}�W���Y���R��d1����u������/���!����kD��N��U���0�1�6�&�l�}�Wϻ�Ӗ��P��d��Uʓ�
�
� �c�`�-�W��
����\��h����� �&�2�0��-��������9��G��U���<�;�1�!�'�n�(���O�ד�O�=N��U���3�
�a�
�e�a�W���&����P9��T��]���<�;�1�4��2�����ԓ� U�N�����0�}�8�
��(�B���	���9F�?��;����d�3�
�n��E��Y���D��F�����}�g�d�3��e�(��Y�ƿ�T�������!�9�d�
�g�t����Y���9F�?��;����3�
�a��o�K���H�ƻ�V�D�����g�3�
�a��o�W���������T�����d�
�c�|�2�.�W��B���4��P�����:�0�
�
�"�l�Bف�K�����1��*���e�%�u�;�w�0�(�������P��G�U����;�0�
�;�����K����V��h�I����;�0�
�;�����H����U��X�����;�u�4�2�f�<��������U��^�����_�u�u�4�0�l��������9��h_�����l�l�%�u�j�u����&¹��l ��V�*��4�1��;�2���������l��E��F��|�_�u�u�6�:�F�������@9��^_�� ��a�
�f�i�w�}�W���YӴ��T��V�����
�
� �d�`��Eϩ�����A9��Y
�*���3�
�e�l�'�u�^��^���V
��d��U���u�&�9�!�'�e����H�ӓ� ]ǻN�����d�4�9�:�2��(���L����Q��h�I���6�'�,�d�>�;�(��M����R��e��ۊ�9�
�;�&�e�4����O�ԓ� O��N��'���0�
�9�
�9�.�E�������
T��N�U���u�u�u��9�8�(���&����l ��X�*��"�0�u�:��2��������P��h�E���u�d�|�0�$�}�W���Y����V
��Z�*���d�m�
�f�]�}�W����ד�_
��Y��G���-�<�
� �f�n�(��E����R��1�����0�
�
�d�%�:�D��Y����P��N1�����<�
� �d�e��E��Y����R��1�����0�
�
� �����Lǹ��Z�<�����4�9�:�0���(���H����CU��Y
�����
�
�:�
��(�F��&���9F�<�����4�9�:�0�����IĹ��Z���B���
�e�d�%�w�3�W���&�ד�F9�� 1��\�ߊu�u�4�2�f�<��������U��Y�����h�w�w�"�2�}����
����9��P1�C���u�%�6�;�#�1�D��Y����D��d��Uʇ�;�0�
�9��3��������S��N�U��u�=�;�}��8����M����lR��N�����:�&�
�#��t����Y���9F�<�����4�9�:�0��(�F��&���F��V ��G���9�:�0�
�����Hù����<�����4�9�:�0�����LŹ��]ǻN�����d�4�9�/�%�.�F���&����l��S��D���=�;�}�4�����@˹��[��G1�����9�`�
�|�2�.�W��B���4��P�����/�'�&�g�1��G���	���N��Y	��*���
�;�&�f�1��G���	�ƴ�AF��h�����#�
�|�_�w�}����H����l��X��*���3�
�d�l�'�}�J�ԜY���F��V��D���
�e�f�%�w�5��������W_��^_�� ��c�
�g�e�w�}�F�������9F�N��U���
�8�f�
�"�l�Bށ�J���F��Y	��*���
�0�:�
�����I˹��Z�=N��U���u�
�m�<�1��A���	�ƻ�V�X�����f�<�3�
�a�e����P���A�R��U���u�u�u�&�;�)��������V��UךU���4�2�d�4�;�'����J����W��h�I���d�u�=�;��<�(���&����U��N�����:�&�
�#�c�m�W�������l�N�����
�9�
�0�8��(���J����CT�
N��Wʢ�0�u�%��$�1�(ށ�����R������!�9�f�e�w�1����[���F��Y	��*���
�0�:�
��(�D��&���F�N�����%��&�9������K�����T�����f�e�u�9�2��U�ԜY�ƞ�]��h��*���:�
� �d�d��E��Y۴��T��V�����
�
� �d�b��EϦ�Ӈ��P	��C1��D��n�u�u��9�8�(���&����_��G\��Hʦ�1�9�2�6�!�>��������A��CF�����0�}�4�
��(�F��&���G	��Y�����;�<�;�1�p�z�QϪ�	����U��V�����d�d�1�"�#�}�^���P���F��Y	��*���
� �d�a��o�K�������T��A�����=�3�
�<�?�u��������R��hX�� ��f�%�|�!��3����Q����T��I�U���8�
�c�3��m�N���Q�����Y��E���|�n�u�u��3�݁�����V��h��D���
�g�i�u�f�}����Q����VT��h]�� ��a�
�g�h�%��F���&����l�������w�_�u�u�6�:�E�������@9��^_�� ��c�
�f�i�w�}�W���YӴ��T��V�����
�
� �d�b��Eϩ�����A9��Y
�*���3�
�e�f�'�u�^��^���V
��d��U���u�'�#�
�"�l�Eށ�K���F��Y	��*���
�;�&�d�>�;�(��I����[�N��U����;�0�
�;���������R��N�����:�
�:�1�f�4����L�ԓ�N��S��D���0�&�u�u�w�}�WϬ�¹��lW��1��N���u��;�0��1�(���
�ד�\��1��*��c�%�u�h��<��������]��1��*���
�l�d�-�%�<�(���
����9��d��Uʇ�;�0�
�9��3��������l ��Y�*��i�u��;�2���������l��B1�Dڊ�f�-�'�4��2����¹��l�N�����
�9�
�;�$�n����I�ד�F�L�U���;�}�
�0�"�)���&����W��S�����;�!�9�g�d�}����[����F�e��؊�9�
�;�&�c�;�(��I����[�L�����}�
�0� �#�n����M����F��h�����#�
�|�0�$�}�G��Y����R��1�����0�
� �d�g��E��Y���D��F�����
�
�
� �f�d�(��DӔ��l ��[�*��u�9�0�w�u�W�W���T�ƭ�l��RN�����u�'�6�&�y�p�}���Y����\��V�����'�6�o�%�8�8�ǿ�&���R��^	������
�!�e�1�0�F���Y����V��=N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�e�����@���G��d��U���u�u�u�4��2���Y����\��h�����n�u�u�u�w�8����Y���F�N�����;�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�<�9�w�.����	����@�CךU���%�<�9�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E�ߊu�u�0�<�]�}�W���Y�����F��*���&�
�:�<��}�W���
����O��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�~�)����Y���F�N�����9�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����W
��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h�����&�<�;�%�8�8����T�����E�����&�2�
�'�4�g��������C9��N��*���
�&�$���)�G�������9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����_�N�����u�u�u�u�w�}��������[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�0�3�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������_��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��^�����2�
�'�6�m�-����
ۇ��@��CB��*ڊ�0�
�9�=��-��������TJ��h_�����4�
�%�#�3�4�(���UӖ��l6��^�����9�
�;�&�0�}�(ځ�����G��G1�����
�<�|�u�w�?����Y���F�N��U���%�&�2�7�3�l�N��Y�μ�9��Q1�����%�#�1�<��4�W���	����@��X	��*���:�u�%�g��/����	����l��D��Hʴ�
�:�&�
�8�4�(�������lW��R�����%�#�1�<��4�W���	����@��X	��*���:�u�%�e�%�;��������E
��^ �����u�%�6�;�#�1����I�ƣ�N��h�����u�%�6�;�#�1����I����F�R �����0�&�_�_�w�}�ZϿ�&����Q��\����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h-�����_�u�u�0�>�W�W���Y���F�N��*���
�1�
�g�w�`�_�������l
��h_��U����
�&�}�w�2����O����F�R �����0�&�_�_�w�}�ZϿ�&����Q��Z����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h-�����_�u�u�0�>�W�W���Y���F�N��*���
�1�
�a�w�`�_�������l
��h_��U����
�&�}�w�2����N����F�R �����0�&�_�_�w�}�ZϿ�&����Q��W����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h-�����_�u�u�0�>�W�W���Y���F�N��*���
�1�
�l�w�`�_�������l
��h_��U����
�&�}�w�2����A����F�R �����0�&�_�_�w�}�ZϿ�&����Q��_�U���<�;�%�:�2�.�W��Y����C9��P1����g�
�&�<�9�-����Y����V��V��&���8�_�u�u�2�4�}���Y���F�N�����<�
�1�
�f�j�K�������]��[��D��4�
��3�:�l��������]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��D���4�&�2�u�%�>���T���F��h��*���
�d�`�4�$�:�(�������A	��D�����
�&�|�u�w�?����Y���F�N��U���%�&�2�7�3�o�D���D�έ�l��D��ۊ�u�u�%���.�_�������T�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����a�u�&�<�9�-����
���9F������7�1�g�a��.����	����	F��X��´�
��3�8�]�}�W������F�N��U���u�4�
�<��9�(��J�����T�����d�d�h�4������Jӂ��]��G����u�;�u�'�4�.�L�ԶY���F��h��*���
�d�e�4�$�:�W�������K��N�����<�
�1�
�f�m��������\������}�%��
�$�t�W�������9F�N��U���u�u�u�%�$�:����K����[�V�����
�#�
�u�w�-�4���
����W	��C��\��u�u�0�1�'�2����s���F������7�1�g�`�w�.����	����@�CךU���%�&�2�7�3�o�Bׁ�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������^�
N�����;�!�9�d�f�`����*����S��X�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�e�}����Ӗ��P��N����u�%�&�2�5�9�E�������]9��X��U���6�&�}�%������Y����V��=N��U���u�u�u�u�w�-��������U�
N�����;�!�9�d�f�`����*����_��X����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�c�}����Ӗ��P��N����u�%�&�2�5�9�E�������]9��X��U���6�&�}�%������Y����V��=N��U���u�u�u�u�w�-��������S�
N�����;�!�9�d�f�`����*����W��S�����e�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��k�W�������A	��D�X�ߊu�u�%�&�0�?���N����Z��G��U���'�6�&�}�'��(���P�����^ ךU���u�u�u�u�w�}��������lT��R��]���6�;�!�9�f�l�JϿ�&����@�N�����u�d�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��F���
������T��[���_�u�u�%�$�:����J�ӓ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��[��H���%�6�;�!�;�l�F������l ��_����!�u�g�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h]�U��}�%�6�;�#�1�F��DӇ��p5��D��Fʱ�"�!�u�f�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����J�ƭ�@�������{�x�_�u�w�-�������� _��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��F���h�}�%�6�9�)����H����C9��h��]���1�"�!�u�b�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lU��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*���u�h�}�%�4�3����H�����t=�����c�1�"�!�w�k�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����������^	�����0�&�u�x�w�}��������W9��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��i�u�4�
��;�������\F��S�����;�!�9�d�f�f�W�������A	��D����u�x�u�%�$�:����J����@��YN�����&�u�x�u�w�<�(���&���� Q��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��F���i�u�4�
�8�.�(���&���R��d1����u�:�;�:�f�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����g�i�u�4��2����¹��F��h-�����d�u�:�;�8�l�^��Y����]��E����_�u�u�x�w�-��������R��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��Z�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����a�a�i�u�6�����&����F�V��&���8�d�u�:�9�2�F���B����������n�_�u�u�z�}��������lR�������%�:�0�&�w�p�W�������T9��S1�B���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�a�b�i�w�<�(���
����9��
N��*���3�8�d�u�8�3���P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��N�����u�'�6�&�y�p�}���Y����Z��S
��A���&�2�
�'�4�g��������C9��V��U���&�2�6�0��	��������F��1�����%�4�4�
�;�t�W�������9F�N��U���u�u�u�%�$�:����L���N��G1�����9�2�6�d�j�-�G�������[��G1�����;�u�:�}��-��������Z��S�����2�6�0�
��.�F������R�������!�9�2�6�g�`��������O�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��4�&�2�u�%�>���T���F��h��*���
�f�4�&�0�����CӖ��P�������!�u�%�&�0�>����-����l ��h^����'�3�8�-�6�����Y����V��=N��U���u�u�u�u�w�-�������� F�F�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�f�/��������E
��UךU���;�u�'�6�$�f�}���Y���R��^	�����g�4�&�2�w�/����W���F�V�����1�
�g�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�g��'�:��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����T�
N�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u����������E
��UךU���;�u�'�6�$�f�}���Y���R��^	�����`�4�&�2�w�/����W���F�V�����1�
�`�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��Yʥ�`�'�3�7�#��������F��P��U���u�u�u�u�w�}��������W9��R��]���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(���&����l��A��\�ߊu�u�;�u�%�>���s���K�V�����&�$��
�#�m����@Ӈ��Z��G�����u�x�u�u�6�����
����g9��^�����
�&�<�;�'�2�W�������@N��h��*���
�g�|�u�w�?����Y���F��QN�����2�7�1�g�d�}����s���F�N�����<�
�&�$����������Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����9��Z1�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���
�&�$���)�F�������R��P �����&�{�x�_�w�}��������B9��h��D���8�d�
�&�>�3����Y�Ƽ�\��DF��*���
�1�
�a�~�}�Wϼ���ƹF�N�����%�&�2�7�3�o�B������F�N��U���4�
�<�
�$�,�$����ד�@��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����
����g9��_�����e�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�<�
�$�,�$����ԓ�@��N�����u�'�6�&�y�p�}���Y����Z��D��&���!�g�3�8�f���������PF��G�����4�
�<�
�3��A���Y����V��=N��U���u�3�}�%�$�:����K���G��d��U���u�u�u�4��4�(�������@��h��*��i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϿ�&����P��h=����
�&�
�d�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��h��*��4�&�2�u�%�>���T���F��h��*���$��
�!�d�;���&����T��E��Oʥ�:�0�&�4��4�(���&����9F����ߊu�u�u�u�1�u��������lU��N�����u�u�u�u�w�}��������V��c1��Dي�&�
�g�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�d�
�$��E��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��Dފ�&�
�f�4�$�:�W�������K��N�����<�
�&�$���������� 9��D��*���6�o�%�:�2�.��������W9�� GךU���0�<�_�u�w�}�W���Q����Z��S
��G���!�0�u�u�w�}�W���YӇ��@��T��*���&�d�
�&��n�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�l�(���&���F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�d�
�&��i�����Ƽ�\��D@��X���u�4�
�<��.����&����l ��h_�����2�
�'�6�m�-����
ۇ��@��U
��A��_�u�u�0�>�W�W���Y�ƥ�N��h��*���
�a�|�!�2�}�W���Y���F��G1�����0�
��&�f�����M���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�&�2�6�2��#���Hƹ��^9��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����0�
��&�f�����LӇ��Z��G�����u�x�u�u�6�����
����g9��X�����`�4�&�2��/���	����@��G1�����1�f�l�_�w�}����s���F�^�����<�
�1�
�d�t����Y���F�N��U���&�2�6�0��	���&����S�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�%�$�:����&����GW��Q��D���h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���&�2�6�0��	���&����P��D��ʥ�:�0�&�u�z�}�WϿ�&����P��h=����
�&�
�c�6�.���������T��]���&�2�7�1�d�l�}���Y����]l�N��Uʼ�u�4�
�<��9�(��PӒ��]FǻN��U���u�u�%�&�0�>����-����9��Z1�U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}��������B9��h��B���8�d�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�>����-����9��Z1�U���<�;�%�:�2�.�W��Y����C9��P1������&�d�
�$��@���
����C��T�����&�}�%�&�0�?���K���F��P��U���u�u�<�u�6���������O��_�����u�u�u�u�w�-��������`2��C_�����d�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����Z��D��&���!�m�3�8�f�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��C_�����d�u�&�<�9�-����
���9F������6�0�
��$�l�(���&�ޓ�@��Y1�����u�'�6�&��-��������S�N�����;�u�u�u�w�4�Wǿ�&����Q��Y�U���;�_�u�u�w�}�W���	����l��F1��*���l�3�8�d�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h��*���$��
�!�n�;���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��F1��*���
�&�
�u�$�4�Ϯ�����F�=N��U���&�2�6�0��	��������l��^	�����u�u�'�6�$�u��������lU��=N��U���<�_�u�u�w�}����	����l��h]�U���;�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������B9��h��E���8�d�u�&�>�3�������KǻN�����2�6�0�
��.�E߁�
����l��^	�����u�u�'�6�$�u��������lR��d��Uʷ�2�;�u�u�w�}��������T9��S1�B���=�;�_�u�w�}�W���Y����Z��D��&���!�e�3�8�f�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�m����H�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�
�&�
�w�.����	����@�CךU���%�&�2�6�2��#���K����lW��D�����:�u�u�'�4�.�_���
����W��\����u�0�<�_�w�}�W����έ�l��h��*��b�u�=�;�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�1��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�
�&�
�w�.����	����@�CךU���%�&�2�6�2��#���J����lT��D�����:�u�u�'�4�.�_���
����W��]����u�0�<�_�w�}�W����έ�l��h��*��`�u�=�;�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�1��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�
�&�
�w�.����	����@�CךU���%�&�2�6�2��#���M����lU��D�����:�u�u�'�4�.�_���
����W��Z����u�0�<�_�w�}�W����έ�l��h��*��f�u�=�;�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�1��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�
�&�
�w�.����	����@�CךU���%�&�2�6�2��#���L����lR��D�����:�u�u�'�4�.�_���
����W��[����u�0�<�_�w�}�W����έ�l��h��*��e�u�=�;�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�1��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�
�&�
�w�.����	����@�CךU���%�&�2�6�2��#���O����lS��D�����:�u�u�'�4�.�_���
����W��[����u�0�<�_�w�}�W����έ�l��h��*��m�u�=�;�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�1��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�
�&�
�w�.����	����@�CךU���%�&�2�6�2��#���N����lP��D�����:�u�u�'�4�.�_���
����W��W��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��D��u�=�;�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��F1��*���
�&�
�u�$�4�Ϯ�����F�=N��U���&�2�6�0��	��������l��^	�����u�u�'�6�$�u��������lW��d��Uʷ�2�;�u�u�w�}��������T9��S1�D���=�;�_�u�w�}�W���Y����Z��D��&���!�
�&�
�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h��*���$��
�!��.�(���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����@��d:��ӊ�&�
�u�&�>�3�������KǻN�����2�6�0�
��.�N����ޓ�@��Y1�����u�'�6�&��-��������
S�N�����;�u�u�u�w�4�Wǿ�&����Q��W�U���;�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�8�1����6����A��R����� �9�d�3��h�B���Y���G��Z�����`�b�%�u�8�}��������EW��UךU���:�9�-���)�0�������A9��B�����
�a�c�%�w�`�_���&����A��^�U���u�%�6�;�#�1�F��B�����[1��0���!��0�!�%��(�������U��[�����h�}�9�
�"�o�Bށ�KӞ����T�����d�d�n�u�w�?����¹��lT��1��U��}�8�d�
�"�o�Cف�KӉ��Q��E	��B���8�'�4�
�f�;�(��K����l�N�����0�e�1�8�%�<�(�������T��N�U»�"�<�;�<�����L������
�����
�;�&�g�1��F���	����F�U�����e�1�8�'�6��E���&����l��S�����<�;�<�
��(�D��&����]��R�����;�&�f�3��o�C���P���F��Z�����1�8�'�4�����O����Z������
�0�
�e�a�<�ϰ�����Q��1����`�|�_�u�w�/����@Ĺ��^	��V ��D���
�e�g�%�w�`�_���
����Z��h��D��
�f�4�1�3�1��������9��h��D��
�g�n�u�w�?�����ѓ�V��P�����
�d�d�%�w�`�_���
����Z��R	��L��4�1�1�9�#�9����&ù��U��X�����_�u�u�'�2�:�N؁�H����V��h�I���7�8�'�0�`�9��������l ��^�*��-�'�4�
�8�.�(���&����F�U�����b�<�3�
�f�k����D�ή�^��RW�����'�4�
�
�"�o�Eށ�KӞ����T�����d�d�n�u�w�?�����ߓ�9��h_�D���u�h�}�4�%��(���&�ד�F9��^��Gʺ�u�4�2�g�6�1����&¹��G9��h��D��
�g�n�u�w�?�����ߓ�l ��Y�*��i�u�6�'�.�l��������Q��h����4�2�g�4�;�2����&����Z9��h_�G���|�_�u�u�%�8��������9��R��]���a�3�
�d�g�-�W�������T��h
�����;�<�3�
�f�l����s���Q��E	��ۊ� �g�e�
�e�a�Wǰ�����Q��1��*��`�%�u�'�3�1��������lV��X��D���
�e�e�%�~�W�W�������V9��h��G���
�g�i�u�9�*��������A��^�U���%�;�!�<�1��C���	����F�U�����<�
� �f�e��E��Yۈ��@��U��F���
�e�g�%�w�/��������U��_�����_�u�u�'�2�:�(�������R��N�U»�"�<�;�<�����J¹��	��G1�����
� �f�l��o�L���Yӄ��V��h�� ��e�
�g�i�w�3� �������A��W�U���1�9�!�1�-�/��������l ��_�*��n�u�u�7�:�/����¹��lT��1��U��}�;�0�3�8��(���&����	��X�����
�
�0�
�g�k�L���Yӄ��V��h��G���
�a�m�%�w�`�_�������D9��Q��A���%�u�'�:�2�;����&����S��G\����u�'�0�2���D���&����l��S�� ���'�9�"�f�1��F���	�ƣ�	��E�����3�
�d�c�'�t�}���Y����A��^1��*���f�a�
�g�k�}��������lR��B1�Fӊ�g�:�u�#�%�1� �������S��G�U���7�8�'�0�>�4����H�ޓ�F�F�����9�"�3�
�f�o����Ӊ��A ��@1��*��`�%�|�_�w�}����&����l��E��E��u�8�
�e��(�D��&���K�
�����e�n�_�u�w�p����I����
9��S�����&�<�;�%�8�8����T�����h^��G���4�1�0�&��.����	����	F��X��´�
�<�
�&�&��(���M����lW�������6�0�
��$�l�(���&���R��^	������
�!�`�1�0�F���Y����V��=N��U���u�3�}�4��2��������F�V�����&�$��
�#�k����H���G��d��U���u�u�u�7�1�m�F��&����V��R�����:�&�
�#�c�o�E��Hӂ��]��G�U���u�u�0�&�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���L����lW��N�����u�u�u�u�w�}����I����
9��S�����h�4�
�:�$�����H���W��X����n�u�u�u�w�8����Qۇ��P	��C1�����d�h�4�
�>�����*����R��D��F���!�0�u�u�w�}�W���Yӄ��lV��Z�����0�&�u�h�6�����&����lV�C��U���;�:�e�n�w�}�W�������9F�N��U���u� �
�
�e�d��������[�o6�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�"��(��@������^	�����0�&�u�x�w�}����I����
9��1�����
�'�6�o�'�2��������F��h��*���$��
�!�`�;���P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�l�(���&���F��R ��U���u�u�u�u�5�;�G��Mʹ��F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�7�3�g�l�Cց������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����9��W�����&�<�;�%�8�8����T�����h^��G���6�d�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����ғ�@��B�����2�6�0�
��.�Fف�
����F��h��*���$��
�!�b�;���P�����^ ךU���u�u�3�}��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�C�������F��F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��D܊�&�
�`�|�8�}�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����R�G�����_�u�u�u�w�}�W���&ù��_��R_��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�(�(߁�K�ߓ�VW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h^��G���1�u�&�<�9�-����
���9F���*ڊ�g�l�1�
�$�4��������C��R�����!��&�
�#�(����&����A��\�Yʴ�
�<�
�&�&��(���M����lW�������4�0��'�4�(���A����lR��B�����2�6�0�
��.�Fف�
����F��h��*���$��
�!�b�;���Uӏ��P��V��&���6� �0�d�b�;�(��O����9F����ߊu�u�u�u�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���O����lW��N�����u�u�u�u�w�}����I����
9��R�����!��&�
�#�(����&����A��\�N���u�u�u�0�$�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����ӓ�@��G�����u�u�u�u�w�}�Wϼ��֓�R��S_��Hʼ�
�!��&��)��������9��P1�F��u�u�u�u�2�.��������]��[����h�4�
�<��.����&����l ��h_�\ʡ�0�u�u�u�w�}�W�������lW��1��U��<�
�!��$���������^��Q��C���%�n�u�u�w�}����Y���F�N��U���
�
�g�l�3�}�J���!����k>��o6��-���������/���s���F�R ����_�u�u�;�w�/����B��ƹF�N�����d�a�
�0�w�.����	����@�CךU��� �
�
�g�n�*�F���
����C��T�����&�}�%�6�{�<�(���&����l5��D�*���
�f�u�%�$�:����&����GW��Q��D���4�
�<�
�$�,�$����ӓ�@��GךU���0�<�_�u�w�}�W���Q����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����R��D��F���:�u�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(��PӉ��N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��1����|�|�u�=�9�W�W���Y���F��Q1��D��
�0�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ʈ�U9��\�*���u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǻN�����
�
� �f�a��E��Yے��lW��h��*��a�4�1�!�'�d�(���J����CT�=N��U���'�
�
�d�1��O���	���N��[1�����3�
�m�d�'�}�����Г�F9��]��G��u�u�6�'�.�l����&����l��S�����!�%�
� �f�l�(������^��B1�BҊ�g�n�u�u�4�/��������9��h_�E���u�h�}�8�o�;�(��L����\��Z��Fۊ� �d�f�
�d�f�W�������lW��X��*���d�f�
�g�k�}����&����U��G\��ʡ�%�b�
� �f�d�(��B�����E��*���f�a�
�g�k�}����H�ޓ�V��W����!�%�l�
�"�n�Dց�K��ƹF��V��*���g�l�
�g�k�}����H�Փ�F9��^��Fʴ�1�!�%�b��(�E��&���9F�
�����;�d�3�
�o��G��Y����w/��x��D���'�2�f�d�l�}�WϺ�����]9��hZ�*��i�u��-��$����K¹��T9��Y�U���1�9�!�1�8�8�(߁�H����_��h�I���1�9�!�1�8�8�(ށ�����9�������!�%�e�3��d�G���P���F��[�����0�
�
�
�"�o�Aׁ�K�����R��*���&�'�2�f�o�}�ϭ�����V��B1�Cي�g�n�u�u�3�1��������9��h_�G���u�h�_�u�w�}�W����ד�_
��Y��G���-�<�
� �f�n�(��������R��Lӊ�d�3�
�l�f�-�_���D����F��D��U���u�u�%�l��l����J����9F�
�����
�;�&�g�1��F���	���l�N��Uʥ�a�
�d�3��m�N���Y����N��E��D���
�e�c�%��t�J���^�Ʃ�@�N��U����;�0�
�;�����L���� V��h����u�0�0�0��3��������R��N�U���u�u�u�%�c��E���&����l��@��U¶�'�,�g�3��o�B���Q���A��N�����u�u�u�u��3�ށ�����V��h��F���
�g�_�u�w�8����&����l ��Y�*��i�u�u�u�w�}�%���¹��_9��R��*���
�
� �d�b��Eϩ�����A��P�*��� �d�a�
�e�m�W���H����_��=N��U���u�
�c�<�1��@���	��ƹF��R�����0�:�
�
�8��F���&����l��S�����c�
�0�
�n�i��������V��R��*ۊ�:�
� �d�n��E��Y����V
��R
�����
�
�:�
��(�E��&���F��Z��F���2�f�b�u�9�}��������A	��Y�����e�`�%�|�]�}�W�������I��D1�����l�f�%�u�j�W�W���Y�ƞ�]��h��*���&�g�<�
�2��N��������E��*���3�
�m�l�'�u�^��^���V
��d��U���u��;�0��1�(�������ZW��R	��L��_�u�u�0�2�8�(�������]	��Q��L���%�u�h�}�2�8��������9��h_�F���u�:�u�%�4�3����H���9F�
�����
�0�:�
��(�E��&���F��^	����� �g�e�
�d�%�ϰ�����A��B1�Eފ�g�n�u�u�3�1��������lU��B1�M܊�f�i�u�u�w�}�Wό�����R
��X ��*ߊ� �f�b�
�e�*��������lW��B1�C܊�g�e�u�u�f�t����Y���F�<�����4�9�/�'�$�i����I�ד�]ǻN�����0�
�0�:�����Oƹ��Z�=N��U���u�4�2�d�6�1����&Ź��lU��1��U���;�}�4�'�����Mƹ��V�
N��R���9�0�_�u�w�}�W����ד�_
��R��*ߊ� �f�c�
�e�W�W�������W9��E�����b�c�%�u�j�W�W���Y�ƞ�]��h��*���&�g�<�3��k�E���Y����N��E��D���3�
�a�a�'�u�^��^���V
��d��U���u��;�0��1�(�������Z9��h_�M���n�u�u�1�;�)��������\��B1�Lߊ�g�i�u�1�;�)��������V��V����4�
�:�&��+�(���s���V��T��*���f�g�
�g�k�}�F������Z*��^1�����:�
�
�0��h�W���	����@��A\��\ʰ�&�u�e�n�w�}����/�ד�F9��1��U��&�1�9�2�4�+����Q����T����*���3�
�a�
�f�}�W���������T�����d�
�e�|�l�}�Wϻ�	����F9�� 1��U��&�1�9�2�4�+����Q����T����*܊� �`�f�%�~�v��������R��X ��*���g��d�|�]�}�W���&����e9��Q��Fۊ�a�i�u�'�0��F���&����CW�N�����u�g�n�u�w�8����	����F9��1��U��<�0�
�
�"�i�@���Q����\��XN�\�ߊu�u�-�
��%��������G��V��*���d�3�
�a�f�-�W��s���F�G1��؊�c�'�2�a�e�}����Q����R��B1�Gۊ�g�e�u�u�f�t����Y���F���*���-� �
�7�8�(��������9��Q��A���%�n�u�u�1�-�6���6����Q��B��#���0�l�
�
�"�o�Eف�K���@��[�����6�:�}�;�>�3�ǿ�&����G9��Z��\��� �&�2�0������HŹ��T9��\��N���u�3�%�������
����V9��[��Lӊ�
� �g�a��n�K���Y���F��h8��G��
� �g�e��n� ���Yے��lQ��Q��@���%�}�|�h�p�z�W������F�N�������!��$�1��������
_��h��G��
�g�_�u�w�%�(�������r��[��*��� �
�l�&�1��B���	�����h�����0�!�'� �$�:����	����@��A\��E���u�;�<�;�3�-�!���&�ד�F9��W��F���_�u�u�-��2��������9��Q��C���%�u�h�&�3�1��������AN��D�����%�6�;�!�;�o�(���Tӓ��Z��SF�����1�
�0�8�b�m�!���&����l��UךU���-�
�:�0�#�/�(��&����lT��1��U��&�1�9�2�4�+����Q����T�������!�9�g�
�~�p��������U��Y��*���8�`�c��1��A���	���9F�N��U���
�:�0�!�%��Gف�&����P��G_��Hʦ�1�9�2�6�!�>����������Y�����9�
�d�'�0�i�A���K���9l�N��Uʳ�%�;�1�
�2�0�B���/����P��h�I���!�
�:�<��8��������VN��P ��]���4�g�d�
�2��G��U���lǻN�����0�8�
�a�����N˹��Z�=N��U���u�
�4�g�f���������9�������0�
�8�a��(�E��&���F�_��U���0�_�u�u�w�}��������U��[����u�u�3�%�/��#�������G��N1�A���3�
�m�a�'�}�JϪ�	����U��X�����g�x�d�1� �)�W���s���U��O#��!���!��9�<�;��Eہ�&����P��G_��Hʧ��a�3�
�o�j���Y����K��z;�����
� �!�%�.�l�C�������R��N�U���
�:�<�
�2�)�Ǭ�
����F��P ��]���
�:�<�
�2�)�ǭ�����U��O#��!���!��9�<�;��Eہ�&����P��G^��_ʦ�2�0�}�-���;�������_��[��Gފ�
� �g�c��l�^��L���9F���*����,� �
�"�)����H�ѓ�l ��V�*��i�u�8�
�n�;�(��H���� T�_�����:�e�n�u�w�;����,����F��B�����d�b��3��e�C���Y����l0��h��G���
�g�_�u�w�%�(���5����G9��[�����g�
�
� �e�j�(��E�ƿ�W9��P�����:�}�0�<�2�(�����ο�W9��P�����:�}�<�;�3�;����,����F��B�����d�b��3��e�C���P����Z��SF����� ���!��1����&����e9��h\�A���|�|�u�b�~�W�W���T�ƫ�C9��hZ�*���4�&�2�u�%�>���T���F��G1��*��
�0�4�&�0�����CӖ��P�������6�0�
��$�l����I�ƭ�l�������7�1�d�l�w�-��������`2��CY�����y�4�
�<��.����&����U��B�����2�6�0�
��.�D������R��^	������
�!�
�$��[Ͽ�&����P��h=�����3�8�a�u�'�.��������l��h��*���u�u�7�2�9�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�8�u��������lW��G�����%�6�;�!�;�:���DӇ��@��T��*���&�b�3�8�a�}����	����@��X	��*���u�%�&�2�4�8�(���
�ԓ�@��N��U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�2�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���ǹ��^9����]���6�;�!�9�0�>�F������T9��R��!���`�3�8�a�w�/�_�������l
��^��U���%�&�2�6�2��#���O����lS�G�����_�u�u�u�w�}�W���&����W��RN�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�0�-����N¹��Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�W�������F9��1��U��%�e�'�3�6�-����&����9F�	��*���a�d�%�u�j�-�F�������l��D�����u�x�u�'��(�C����ƭ�@�������{�x�_�u�w�/�(���M�ѓ�V9��D��*���6�o�%�:�2�.��������V��c1��D���8�e�u�%�4�q��������W9��B�����2�6�0�
��.�@������R��^	������
�!�
�$��[Ͽ�&����P��h=�����3�8�g�u�'�.��������l��h��*���4�
�<�
�$�,�$���ƹ��^9�������6�0�
��$�k����L���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u��<�(���
����T��N�����<�
�&�$���ށ�
������ ��]���&�2�7�1�f�d�^ϱ�Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���}�%�6�;�#�1����H����C9��P1������&�g�3�:�l�W���Q����\��h�����u�u�%�&�0�>����-����l ��h\�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t��������]��[����h�4�
�<��.����&����U��G�����%�6�;�!�;�:���DӇ��@��T��*���&�c�3�8�b�t�^Ϫ���ƹF�N��U���'�
� �a�`�>�W������]��[����_�u�u�u�w�1��ԜY���F�N�����
�b�
�0�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R�����u�2�%�3��j�(��E�Ƽ�9��Q1�����;�&�2�_�w�}��������l��S��*ۊ�0�
�4�
�9�.��ԜY�ƥ�l��t��*��� �!�'�
�`��(���J����CT�
N�����2�6�#�6�8�u����ۏ��P��V��&���6� �0�d�o�i����M�ӓ�O������%��9�
��m����M����]ǻN��9���
�4�0��%�>����H�ד�F9��X��F��u�u�u�u�w�3� ���H¹��lU��1��U���;�}�'�6�9�h����L�֓�N��S��D���0�&�u�u�w�}�Wϰ�����9��h]�@���n�u�u�u�w�4�(���:����`��T����m�a�3�
�c�h����Dӕ��l
��^�����'�'�&�/��4��������
9��h]�@���|�f�|�n�]�}�W�������@��C�����
�b�
� �d�j�(��E��ƹF�N�����9�`�3�
�b�j�������\��X ��*���f�f�
�g�g�}�W��PӃ��VFǻN��U���0��9�a�1��B���	��ƹF��{1��*���0��'�6�"�8�F���M���� R��h�I���!�
�:�<��8����
����WN��h��6���
�!� �!�%��@ށ�&����V��G\��Xʦ�2�0�}�
�6�o�Bف�����U�d��Uʼ�
�!��&��)��������9��h]�C���u�h�_�u�w�}�W���*����l ��[�*��"�0�u�:��2�ځ�����9��^��H��r�u�9�0�]�}�W���Y����V
��h��F��
�f�_�u�w���������\��X�� ��g�
�g�i�w�)�(�������P�������1�<�
�<��/�;���&����T9��G��U���<�;�1�4��2��������]ǻN��9���1�
�0�8�f�m����J�֓�F���*���<�
�0�!�%�(�����θ�CW��Q��F���%�|�~� �$�:����&����l��1����d�|�n�u�w�4�(���¹��l4��P�����:�'�0�g�1��@���	���l�N��Uʴ�
�:�&�
�!�o�Gϩ�����V
��Z�����b�d�%�}�~�`�P���Y����l�N��Uʦ�9�!�%�
�"�n�Fہ�J���F�N��*����g��!�e�o����N�֓�F���*���<�
�0�!�%�/����Q����V��Z��EҊ� �f�f�
�c�q�E���s�����O=�����
�e�
� �d�n�(��E�ƿ�W9��P�����:�}�;�<�9�9����)����W9��h��\��� �&�2�0������H����a��R1�����0�6�
�
�"�n�Eف�J����F�^��D���
�e�
�g�k�}�F������@��R
�����f�
� �m�b�-�^��
����WN��h�����#�
�|�u�;�8�U���s���Z��1��*��
�g�i�u�f�}����Q����V��Z��Fي� �l�d�%�~�c�����έ�l��D�����e�|�0�&�w�m�L���Yӏ��CU��Y�����c�l�%�u�j�u����&����^��G\�����%�6�;�!�;�l�F��Y����P��h��G��
�g�i�u�f�}����Q����R��Q��@���%�u�u�%�4�3����K���V
��L�N���u�<�8�
�"�k�N���Y���D��_��]���;�1�!�%�o����@����X��^	��´�
�:�&�
�!�l�G�������V�=N��U���2��d�3��l�(��E�ƨ�R��P ��*���a�c�%�n�w�}����&����lR��h�I���
�&�<�;�1��O܁�H���F��Y��D���
�g�
�f�k�}����/�ד�F9��1��]��1�"�!�u�d�f�W�������U��Y��D��u�8�
�f�1��Nށ�K���W��X����n�u�u�9��(�F��&���F��G1�*���d�a�
�g�f�p�FϺ�����O��=N��U���9�
�
�a���(���������^	�����0�&�u�x�w�}����&����V9��V
�����
�&�<�;�'�2�W�������@N��h��*���$��
�!�`�;���UӇ��@��T��*���&�d�
�&��e�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������D�����
��&�d��.�(��PӒ��]FǻN��U���u�u�!�e�c�h��������@��S�����;�!�9�c��u�W���Y����G	�UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	���&����P����ߊu�u�u�u�w�}����M�ӓ�lV��S
����i�u�%�6�9�)���&����F��S�����|�_�u�u�w�}����s���F�N�����
�a�
�
��9����I���>��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�9�
��i�(���&����V�������%�:�0�&�w�p�W�������R��R1�����0�&�
�&�>�3����Y�Ƽ�\��DF����`�'�2�a�b�q��������V��c1��Dӊ�&�
�m�u�'�.��������l��1����|�u�u�7�0�3�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��M���8�d�|�u�?�3�}���Y���F�[��*��
�
�
�1�%�.�F��Y����V��E��A���}�u�u�u�8�3���B���F������}�%�6�;�#�1����H����C9��P1������&�d�
�$��O�������9F�N��U���u�!�e�a�b�8�G�������F������!�9�c�
��}�W�������V�=N��U���u�9�0�_�w�}�W���Y�Ơ�lV��[��*ڊ�1�'�&�d�k�}�/���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*ڊ�a�
�
�
�2�}����Ӗ��P��N����u�!�e�a�b�8�G���I����Z��G��U���'�6�&�}�'�>�[Ͽ�&����P��h=����
�&�
�c�w�-��������`2��C_�����d�|�u�u�5�:����Y�����F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�/�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���@����lW��G�����u�u�u�u�w�}�Wϲ�&ù��9��1��E��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����&����V9��T�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*ڊ�a�
�
�
�2�}����Ӗ��P��N����u�!�e�a�b�8�G���H����Z��G��U���'�6�&�}�'�>�[Ͽ�&����P��h=����
�&�
�m�w�-��������`2��C_�����d�|�u�u�5�:����Y�����F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�/�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���A����lW��G�����u�u�u�u�w�}�Wϲ�&ù��9��1��D��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}����&����V9��T�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B���F��h^��Aߊ�
�
�d�i�w�0�(��&����U��GZ����u�x�9�
��i�(���&����R��P �����&�{�x�_�w�}����M�ӓ�lV��R_�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�f�����N���F��P��U���u�u�<�u��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�Fׁ�
����O����ߊu�u�u�u�w�}����M�ӓ�lV��R_��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�)�G��L����l��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��C1��A���0�d�4�1�2�.�W�������A	��D�X�ߊu�u�!�e�c�h��������@��V�����'�6�o�%�8�8�ǿ�&����P��h=����
�&�
�c�w�-��������`2��C_�����d�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�5��ԜY���F�N��*ڊ�a�
�
�
�3�/���E�ƭ�l��D�����d�g�x�d�3�*����P���F�N�����}�4�
�:�$�����&���R��^	������
�!�b�1�0�F���Y����l�N��U���u�9�
�
�c��(ށ�����@V�
N��*���&�
�#�a�g�o�Z������\F��d��U���u�0�&�u�w�}�W���Y����G9��Z�����4�1�0�&�w�`�U���B���F���U���u�u�u�0�3�-����
��ƓF�C�����a�`�0�d�6�9����Y����T��E�����x�_�u�u�#�m�C����ד�W��D�����2�
�'�6�m�-����
ے��lW��h��*��m�u�%�&�0�>����-����
9��Z1�Yʴ�
�<�
�&�&��(���A����lW��=N��U���<�_�u�u�w�}��������]��[����h�4�
�<��.����&����l ��h_�\ʡ�0�u�u�u�w�}�W�������R��R1�����0�&�u�h�#�-�F�������S��N�Dʱ�"�!�u�|�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��L���8�d�|�u�?�3�}���Y���F�[��*��
�
�
�1�%�.�F��Y����\��h��A��g�x�d�1� �)�W���s���F�R��U���u�u�u�u�w�1�(߁�Mƹ��9��S�����h�w��n�w�}�W�������U]�N�����%�:�0�&�]�W�W���Tӊ��9��1��D���e�4�&�2�w�/����W���F�[��*��
�
�
�0��.����	����	F��X��´�
�0�u�%�$�:����&����GW��Q��D���4�
�<�
�$�,�$����ߓ�@��GךU���0�<�_�u�w�}�W���Q����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����Q��D��C���:�u�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(��P����[��=N��U���u�u�u�!�g�i�B���H����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�!�e�c�h�������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���Tӊ��9��1��D���d�4�&�2�w�/����W���F�[��*��
�
�
�0��.����	����	F��X��´�
�0�u�%�$�:����&����GW��Q��D���4�
�<�
�$�,�$����ޓ�@�� GךU���0�<�_�u�w�}�W���Q����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����_��D��M���:�u�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(��P����[��=N��U���u�u�u�!�g�i�B���H����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�!�e�c�h�������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�}�Wϲ�&ù��9��1��U��&�1�9�2�4�+����Q����T�������d��
�4�0���������lT��B1�G܊�f�u�u�;�>�3�Ƿ�&����gT��B��D؊� �f�`�
�f�t�}���Y���_��hZ�*���
�0�u�&�>�3�������KǻN�����a�`�0�d� �l��������\������}�%�6�y�6�����
����g9��V�����b�_�u�u�2�4�}���Y���Z �F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��DҊ�&�
�b�|�~�)����Y���F�N�����a�`�0�d� �l�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F���E��`�0�d�"�f�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠu�u�8�;��l����H�ԓ�F���*���<�
�0�!�%�(�����έ�l��D�����e�u�u�;�>�3�Ǯ�+����G9��Q��D���%�|�n�u�w�0����J����P��G\��Hʦ�1�9�2�6�!�>��������V��G1�����9�`�
�|�z�(�����μ�a��[��*���c�f�%�|�l�}�Wϳ�����l ��Y�����h�_�u�u�w�}����&����lP��h����u�<�;�2�f�;�(��&���F�_��U���0�_�u�u�w�}�(�������l ��X����u�u�8�;��;�(��A����[�N��U���8�;��d�1��F���	�ƻ�V�^�����2�f�d�}�~�`�P���Y����l�N��Uʥ��&�9�
��(�F��&����F�Y����
� �f�d��n�K���Y���F��{1��*���0��'�6�"�8�F���M���� R��h����u�&�9�!�'�o����M����O�I�\ʰ�&�u�u�u�w�}��������V9��E�� ���d�`�a�3��i�C���B�����d��D���
�`�g�%�w�`�}���Y���]��R�����a�b�%�u�?�3�_�������l ��Z�*��e�u�u�d�~�8����Y���F��R��Ҋ� �f�e�
�d�W�W�������T��B1�Aފ�f�i�u�u�w�}�WϷ�&����R��d�����0�d�`�a�1��C���	�ƻ�V�D�����d�3�
�a�f�-�_���D����F��D��U���u�u�<�
�#���������F��Y��A���
�a�l�%�l�}�Wϰ����� 9��h]�G���u�h�_�u�w�}�W�������@��C�����
�b�
�
�"�n�Gځ�Hӑ��]F��R�����
� �f�a��o�G���Y�����RNךU���u�u��6��<��������A��[��*���f�d�
�g�]�}�W���*����l ��[�*��i�u�u�u�w�}��������V9��E�� ���d�m�a�3��i�B���Y����N��[1�����'�2�a�e��t�J���^�Ʃ�@�N��U���<�
�!��$���������Q��1��*��l�%�n�u�w�3� ���Hƹ��lU�� 1��U��_�u�u�u�w�8�$���K���� S��h����u�:�
�:�3����@ƹ��V�
N��R���9�0�_�u�w�}�W���*����l ��[�*��_�u�u�0��1�A���&����l��S��U���u�u�<�
�#���������F��Y��A���
�a�`�%�w�5��������CP��Q��A���%�}�|�h�p�z�W������F�N��*����&�
�!�"�)����Aƹ��U��_����u�u�;�"�2�l�(���J����CU�
NךU���u�u��6��<��������A��[��*���f�d�
�g� �8�Wǭ�����T��R	��D��e�u�u�d�~�8����Y���F��{1��*���0��'�6�"�8�F���M���� R��h����u�0��9�o�;�(��A����[�N��U���;�"�0�d��(�D��&����[�������f�3�
�a�b�-�_���D����F��D��U���u�u�<�
�#���������F��Y��A���
�a�l�%�l�}�Wϰ�����l ��Y�*��i�u�u�u�w�}��������G��h[�*��� �g�b�
�e�*��������]��B1�MҊ�g�e�u�u�f�t����Y���F� ��&���3�
�c�f�'�f�W�������_T��B1�Bߊ�f�i�u�u�w�}�Wϸ�	����V9��E��Aڊ�
� �g�`��l� ���Yے��l^��E��A��}�|�h�r�p�}����s���F�Q�����
�0�8�`�f�����O�ד�]ǻN��U���0��9�g��<����&����l��S�����:�<�
�0�#�/�����ο�T�� ��&���
� �g�c��n�[��P��ƹF��R��ي� �g�g�
�d�a�W���Y��� ��h �����'�
�l�
��(�E��&����[����*���`�
� �g�o��E��Y���O��[�����u�u�u�-��2��������9��Q��C���%�n�u�u�9�*�������� R��N�U���u�u�u�3�'�3��������P��h��G��
�d�"�0�w�)���&����V��^��H��r�u�9�0�]�}�W���Y����]	��h����b��3�
�a�o���Y����V��[[�� ��a�
�f�i�w�}�W���Yӈ��`��h��G��
�f�"�0�w�2�(�������P��h�E���u�d�|�0�$�}�W���Y����K��X
�����
�a�
�
�"�o�Bց�H���F��@=��C���
�b�g�%�w�`�}���Y���]��R�F���&�
� �g�`��Fϩ�����A9��Y
�� ��m�
�g�e�w�}�F�������9F�N��U���
�:�0�!�%��N؁�&����P��G\�U���;�"�0�b�1��C���	���l�N��Uʼ�
�!��&��)��������9��Q��A���%�u�=�;��8�(���O¹��lU��1��]���h�r�r�u�;�8�}���Y���Z*��C1�����!� �!�'��j�(ہ�����9��d��Uʻ�"�0�m�3��h�F���Y���F�N�����!��&�
�#�(����&����9��h]�A���u�=�;�}�2����&����R��G\��\��r�r�u�9�2�W�W���Y�ƥ�l��t��*��� �!�'�
�`��(���J����CW��N�����0�l�3�
�`�h����D���F�N��#���
�d�'�2�c�k�W����ο�_9��G[�����c�a�%�}�~�`�P���Y����l�N��Uʥ��9�
�c�%�:�C��B�����d�����c�f�%�u�j�W�W���Y�ƪ�C9��S�����`�c��3��k�O���Y����N��[1�����'�2�a�l��t�J���^�Ʃ�@�N��U���3�%�;�1��8���H����F9�� _��G�ߊu�u�0�&�0�?��������
S��N�U���4�g�d�
�"�l�@݁�J����W	��C��B��u�u�;�"�>�3����&���� Q��G]��Hʥ��9�
�e�1��D���	������Y��G���_�u�u�0�$�:����J���� V��h�I���
�4�g�`��(�D��&���F��@ ��U��n�u�u�;� �4����&ǹ��lU��1��U��%��9�
�d�;�(��O���� W��X����|�_�u�u�8�����&����V��G\��H���0�&�2�7�#�o����J�ޓ� F�������!�d�
�:��(�E��&���9F������d�3�
�b�g�-�W��Q����G��1����l�u�'�<�:�n����M����l�N��*���1�
� �g�f��E��Yۉ��P	��h��G��
�g�:�u�%�>��������V��G�U���:�
�:�1��(�D��&���F��R����
� �f�m��o��������CS��Q��A���%�|�_�u�w�/����M���� S��h�I���&�9�!�%�`�;�(��L����\��Z��Eڊ� �f�d�
�e�f�W�������]��Q��@���%�u�h�}�%�>��������
S��N��U���6�;�a�3��h�N���P���F��h�����<�
� �d�d��E��Yے��lP��Q��E���%�u�;�u�2�n����I�ד�O��N�����:�1�d�<�1��B���	���N��G1�*���d�b�
�g�6�9����&����Q��G\����u�'�6�;�n��F���&����l��S�����c�
� �d�e��EϿ�Ӕ��9��hW�*��n�u�u�:��2��������P��h�I���!�%�g�
�"�l�@ف�KӇ����h��D��
�g�n�u�w�2�(�������P��h�I���&�9�!�%�e�;�(��M����\��R�����
�0�
�e�`�f�W�������_	��1��*��c�%�u�h��/����&�ד�F9��[��Gʴ�1�!�%�b��(�E��&���9F������"�g�3�
�c�j����D�ή�^��R1��*���g�`�
�g�6�9����NĹ��lT��1��\�ߊu�u�#�'�;�*�D���&����l��S�����'�0�<�
�"�n�Eځ�KӇ����hW�����d�d�%�|�]�}�W�������lR��B1�Dߊ�g�i�u�7�:�/����&���� V��G\�����8�
�m�3��n�G���P���F��R����� �g�d�
�e�a�WǼ�����l��B1�Eߊ�g�4�1�!�'�n�(���K����CT�=d��U���u�
�
�0��1����	����l��D�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��Q1�����4�
�9�
�9�.����
����C��T�����&�}�
�
�2�����&����_�G1�����4�%�4�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*ڊ�0�
�9�=��-����PӒ��]FǻN��U���u�u�
�
�2�����&����_��Y1����u�
�
�0��1����	����l�N��Uʰ�&�u�u�u�w�}�W���	�֓�V ��[��*���#�1�<�
�>�}�JϮ�I����l��_�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l��h�����;�&�2�4�$�:�W�������K��N�����'�3�4�%�6�4�(���&����T��E��Oʥ�:�0�&�%�g�/����	���C9��E�����4�%�0�y�'�m��������l��A�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�g�/����	����C9��SG�����u�u�u�u�w�}�WϮ�I����l��_�����2�i�u�
��8�(�����ƹF�N�����_�u�u�u�w�}�W���&����R
��V1��*���u�h�%�e�%�;��������T]ǻN��U���;�u�3�u�w�}����	����@��=N��U���`��6�:�w�`����
����V9��E�� ���d�m�6�&��8�(��@��ƹF�N��Dߊ�0�!�'�4��1�W�������A	��D�X�ߊu�u�
�`��>����	����l��^	�����u�u�'�6�$�u����UӇ��@��T��*���&�g�
�&��d�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�e�1�0�F���PӒ��]FǻN��U���u�u�
�`��>����	����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�
�`��>����	����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lW��R�����%�#�1�<��4�W�������A	��D�X�ߊu�u�
�
�2�����	����l��D�����2�
�'�6�m�-����
ۖ��l��h��*���#�1�u�
��8�(���&����_��E�����u�0�<�_�w�}�W�������C9��Y�����6�d�h�%�f�/��������E
��N�����u�u�u�u�w�}��������R��G1�����
�<�u�h�'�l��������C9��SUךU���u�u�9�0�]�}�W���Y���C9��E�����4�
�9�
�9�.���Y����A��Z�����9�
�'�2�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ƽ�9��Q1�����
�<�u�&�>�3�������KǻN��*ۊ�0�
�4�
�9�.����
����C��T�����&�}�
�
�2����	�ד�V ��V�����u�
�
�0��<�(������F�U�����u�u�u�<�w�u��������\��h_��U���
�0�
�4��-����PӒ��]FǻN��U���u�u�
�
�2���������Z�G1�����8�-�_�u�w�}�W������F�N��Uʥ�d�'�3�8�/�4�(���Y����lW��R�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&����A��h�����<�
�<�u�$�4�Ϯ�����F�=N��U���
�0�<�1�6���������l��^	�����u�u�'�6�$�u�(݁�����l��A��U���
�0�<�1�6��������F�U�����u�u�u�<�w�u��������\��h_��U���
�0�<�1�6�����Y����l�N��U���u�%�g��%�2�(�������]9��PN�U���
�0�<�1�6����Y���F��[�����u�u�u�u�w��(�������C9��S1��*���u�h�%�g��/����	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�
�
�0�>�9��������l*��G1�����c�f�%�u�j�W�W���Y�Ƽ�9��E��*���&�2�"�0�w�)���O���� P��h�E���u�d�|�0�$�}�W���Y����F ��h_�L���n�_�u�u�z�-�E�������Z��^	�����;�%�:�0�$�}�Z���YӖ��l6��^�����<�
�&�<�9�-����Y����V��G1��%���:�y�%�g��/�������C9��g�����%�#�1�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	�ԓ�V��S1��*���|�u�=�;�]�}�W���Y���C9��g�����;�&�2�i�w��(�������F�N�����u�u�u�u�w�}�WϮ�K����Z	��^ �����h�%�g��%�2�(������F�N��ʼ�n�_�u�u�9�}����
��ƓF�G1�����g�d�%�u�j�W�W���Y�ƭ�l��D��������u�?�3�_�������T9��Y��\��r�r�u�9�2�W�W���Y�ƭ�l��D�����e�_�u�u��e�ށ����� 9��R��]���'�
�
� �d�k�(������R��1�����0�
�
� �d�j�(��B�����1��*���f�l�
�g�k�}���� �ԓ�F9��[��Gʴ�1��;�0��1�(���
�Г�F9��[��G��u�u�%�f�����M����Z������0�
�e�b�6�9��������V��]�N���u�%�f�3��j�O���Y���F�N�����:�&�
�#�o�n�1���������R	��*���
�m�l�e�w�}�F�������9F�N��U���6�;�!�9�f��L���YӖ��9��h��F��
�g�i�u��3�݁�����V��h��F��
�g�4�1�#�-�N܁�����9��UךU���
�d�<�
�"�n�@ׁ�K���4��P�����:�0�
�
�"�n�B߁�KӇ����hW�����g�f�%�|�]�}�W���Y����r9��Z��*���u�h�&�1�;�:��������A��M�����1�9�
�
�c��(߁�����V��Y�Y��|�_�_�u�w�p����8����Z��R1�����9�u�&�<�9�-����
���9F���*���<�<�2�0�g�<�(���&����T��E��Oʥ�:�0�&�4��8�W���
����@��d:�����3�8�d�|�w�}�������F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�n�t�W������F�N��Uʥ�a��!�8�9��(߁�	����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�
�
��4�����֓�C9��SN�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���C9��v1�����
�
�u�h�4��9���8����A��\��*ۊ�0�
�g�a�]�}�W��Y����r9��Z��*���
�%�#�1�6�.��������@H�d��Uʥ�a��!�8�9��(ށ�	����l��^	�����u�u�'�6�$�u����UӇ��@��T��*���&�g�
�&��d�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�e�1�0�F���PӒ��]FǻN��U���u�u�
�
��4�����ד�C9��SN�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�'�i�6�������V9��V�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�0�
�0�6�<�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�L����l��V1��*���
�;�&�2�6�.���������T��]���
�0�
�0�6�<�(���UӖ��l��h�����
�9�
�'�0�W�W�������F�N�����}�%�6�;�#�1����H����lS��R�����4�
�9�|�w�5��ԜY���F�N��@���3�7�!�
�'�+����&����[��h[�����0�4�4�
�;�f�W���Y����_��=N��U���u�u�u�
��8�(�������E
��^ �����h�%�`�'�1�?����	����l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��8�(�������@��V�����'�6�&�{�z�W�W���&ƹ��U9��C�����2�4�&�2��/���	����@��h[�����0�4�u�
��8�(�������TJ��h[�����0�4�4�
�;�t�W�������9F�N��U���}�4�
�:�$�����&���C9��E�����
�%�#�1�~�)����Y���F�N��*ߊ�0�
�0�4�>�����DӖ��l��h���ߊu�u�u�u�;�8�}���Y���F�G1�����7�!�
�;�$�:�K���&ƹ��U9��C�����_�u�u�u�w�3�W���Y����������n�_�u�u�w�}�(ف�&����]��h^��Hʦ�1�9�2�6�!�>����������Y�����
�a�
�
��m�[��P��ƓF�C��*܊�
�<�<�2�2�m�����ƭ�@�������{�x�_�u�w��(�������l��h�����4�&�2�
�%�>�MϮ�������T����<�
�&�$����������
OǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���Kù��^9��G�����u�u�u�u�w�}�WϮ�O����Z��P1��E���
�9�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��C�����
�
�%�#�3�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠu�u�%�c��)����&����[��C1��A���0�d�$�n�]�}�W��	�Г�l��^ �����4�
�9�u�$�4�Ϯ�����F�=N��U���
�
�<�<�0�8�F���&����R��P �����o�%�:�0�$�<�(���Y����Z��D��&���!�e�3�8�f�t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��N���Y����l�N��U���u�%�c��#�0����&¹��l��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u���(�������lW��G1����u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��ƓF�N�������8�;���W��
����\��h�����'�&�/�}�>�3�ǲ�&ù��9��1��\��|�n�_�u�w�p�W���&����^��h��*���#�1�4�&�0�}����
���l�N��M����8�;�
����������Z��G��U���'�6�&�}�'�>�[Ͽ�&����P��h=����
�&�
�l�]�}�W������F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�e�3�8�f�t�^Ϫ���ƹF�N��U���
�
�
�<�>�:��������WF������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�%�m��	����&����R��[
��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s�����h-�����2�0�d�i�w�)�G��L����l��=d��U���u�
�
�
�>�4����H����E
��V�����'�6�&�{�z�W�W���&˹��g��Y	��*ۊ�%�#�1�4�$�:�(�������A	��D�����y�4�
�<��.����&����l ��h_����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GT��Q��D���|�!�0�u�w�}�W���Y����l^��h:�����0�d�4�
�;�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�G1��6���8�;�
�
��-����E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�-�Nځ�H����W��h�I����;�0�
�;�����&����lW��1��U���'�#�
� �n�l����s���C9��h�� ��c�
�g�i�w�����&����I��D1�����c�a�%�u�%�/����&����l��d��Uʥ�l�
�d�3��l�B���Y���G��]�����d�b�%�u�%�����&����I��D1�����e�b�%�|�]�}�W���O����F9��V��G��u�!�%�d�b�;�(��I����\��V ��D���9�/�'�&�1��A���	����F�G1�*���3�
�e�f�'�}�J�������l ��^�*��4�1��;�2���������9��h_�B���|�_�u�u��e����&����l��S�����f�
� �d�d��EϿ�Ӵ��T��V�����&�3�
�c�a�-�^�ԜY�Ƽ�a��[��A���!�3�
�f�o�-�W��Q����R��Q��F���%�u�:�u�'�>�����ד�]ǻN��*��� �!�g�3��h�(��E����R��hX�� ��f�%�u�;�w�0�(��&����W��G�U���%��&�9�����A˹��Z�D�����6�#�6�:��8��������]��C��A���
�d�d�%�~�h�^��Y����l4��B��B���
�c�
�d�k�}��������E��X�����0� �&�2�2�u����A����S��G]��@���n�u�u�%��.����&���� R��G\��H���4�
�
� �f�d�(������^��1��*��a�%�|�_�w�}�(���K����^��Q��G���%�u�h�_�w�}�W���	����@��A_��D����"�0�u�5�0��������U��\�����|�h�r�r�w�1��ԜY���F��a��*���'�2�f�l�l�}�WϮ�/����P��B1�Dߊ�f�i�u�u�w�}�WϮ�/����9��O1��*��g�%�u�=�9�u��������U��_�����|�h�r�r�w�1��ԜY���F��[1�����3�
�d�g�'�f�W���	����9��h��D��
�f�i�u�w�}�W�������W��R	��M���"�0�u�&�;�)��������
T��G��U��|�0�&�u�w�}�W���
����^��h��D��
�f�_�u�w�����H����S��h�I���u�u�u�u�6�����&����l^��^����u� �1�'�;�*�E���&����l��G��U��|�0�&�u�w�}�W���	����9��h��*��a�_�u�u��<�E��H����l ��_�*��i�u�u�u�w�}��������_��hY��3����"�0�u�5�0��������U��X�����|�h�r�r�w�1��ԜY���F��a��*���3�
�e�b�'�f�W���	����9��1�����
�f�g�%�w�`�}���Y���R��X ��*���g�b����}����Q����A��^1��*���f�a�
�g�g�}�W��PӃ��VFǻN��U���
�4�g�`��(�D��&����F�G1��؊�f�8�-�3��i�B���Y���F�N�����:�&�
�#�c�j�1���Y����N��Z�����<�
� �g�`��E��Y���O��[�����u�u�u�
�6�o�D߁�����R��N�����9�
�b�3��o�O���Y����K��R��*��
�
� �g�`��D�ԜY�Ƽ�e��h\�����g�m�%�u�j�.��������V��EF�����}�;�<�;�3�.��������V��EF�����}�
�4�g�e����@˹��F�D�����e�u�4�
�8�.�(���L����vO�N�\��u�u�%��;��N���&����l��S��*���g�g�
� �e�d�(��J�ƨ�D��_�N���u�%��9���N���&����l��S��U���u�u�4�
�8�.�(���K����V��N����� �1�'�9� �n����H�֓�N��S��D���0�&�u�u�w�}�WϮ�/����W��B1�A݊�g�_�u�u��<�E�������T��N�U���u�u�u�!�'�o�(���H����CW��_��]���
�
� �d�d��E��Y���O��[�����u�u�u�
��(�F��&����F�G1��؊�e�3�
�f�e�-�W��
����\��h����� �&�2�0������Kʹ��lT��1��\��� �&�2�0��0�(�������^��G����u�
�4�g�d�o�(���J����CU�
NךU���u�u�%�6�9�)���&����V�������;�0�3�:�����Jʹ��V�
N��R���9�0�_�u�w�}�W����ԓ� 9��h]�C���n�u�u�%��1�(܁�����9��R�����9�2�6�#�4�2�_���������V��G���
�g�g�%�~�v��������G��_�� ��m�
�d�|�]�}�W����ԓ�9��h\�L���u�h�_�u�w�}�W����ԓ� 9��O1��*��`�%�u�=�9�u��������9��C1��*��l�%�}�|�j�z�P������F�N�����9�
�
� �e�m�(��s���C9��[\��M���
�b�m�%�w�`�}���Y���]��R�����b�a�%�u�?�3�_�������l ��Y�*��e�u�u�d�~�8����Y���F��O�����!�'�
�e�����O˹��l�N��#���
�
� �d�a��D��Y���F���*���3�
�g�m�'�}����Q����G��1��*��m�%�}�|�j�z�P������F�N�����!�%�f�3��i�B���B�����V��@ۊ� �f�a�
�e�a�W���&����P9��T��]���<�;�1�%��1�(�������T��E�����;�1�!�%�n����M����O��N�����9�
�f�3��o�A���Y����G��X	��*���!�'� �&�0�8�_����ԓ�9��P1�B���~� �&�2�2�u����L���� T��h�\�ߊu�u�
�4�e�h�(���J����CU�
NךU���u�u�
�4�e�o�B������� U��h����u� �1�'�;�*�C������� U��h�E���u�d�|�0�$�}�W���Y����l0��1��Gۊ� �f�b�
�d�W�W���&����lS�� 1��*��l�%�u�h�]�}�W���Y����V
��Q��B���%�u�=�;��/����K����Q��h�E���u�d�|�0�$�}�W���Y����V��[Z�� ��f�
�f�_�w�}�(���K�ӓ�F9��W��F��u�u�u�u�w�<�(���
����R�������8�
�
�0��e�E��Y���O��[�����u�u�u�%�4�3����Kǹ��V��d��Uʥ��9�
�
�"����O����Z�=N��U���u�%�6�;�#�1�Eہ�?������YN�����2�
�
�
�"�o�Dׁ�K���F�G�����_�u�u�u�w�����M����lU��UךU���
�4�g�c�1��O���	�����h�����0�!�'� �$�:����&����l_��B1�Lߊ�f�u�u�;�>�3�Ǫ�	����U��\�����n�u�u�%��1�(؁�����9��R�����u�u�u�-��2��������9��Q��C���%�u�=�;��/����&����^��G\��\��r�r�u�9�2�W�W���Y�Ƣ�D5��h��G��
�f�_�u�w�����A����Q��h�I���u�u�u�u�9�*��������T��N�����:�
�:�1��(�E��&���F�_��U���0�_�u�u�w�}��������lT��1��N���u�%��9�����@ƹ��Z�=N��U���u�8�
�g��8�(��Iӑ��]F��Z��F���2�f�m�}�~�`�P���Y����l�N��Uʥ�f�3�
�b�o�-�L���YӖ��R
��D1�*���f�l�
�f�k�}�W���Y����l0��1�D���-�3�
�d�d�-�W����ι�W��[��F���!�3�
�d�`�-�_���D����F��D��U���u�u�%��;��(�������
W��UךU���
�4�g�&�1��E���	���l�N��Uʴ�
�:�&�
�!�e�Gϩ�����^��1����b�}�|�h�p�z�W������F�N��*���&�
�#�m�e�m�G�ԜY�Ƽ�Z*��C1�����:�
�4�!�1��A���	�����h�����0�!�'�'�$�'�_���������{1��*���
�:�%�&�1��A���	���O�=N��U����9�
�:��2��������W��N�U���u�u�u�4��2�����ד���YN�����c�
� �f�a��D��Y���O��[�����u�u�u�8��k�(���J����CW��N�����!�<�
� �d�l�(��E����V
��R
�����
�
� �f�o��DϦ�Ӈ��P	��C1��D��n�u�u�%�9�)�݁�����9��R��]���0�0�
�0�8��(���J����CU��X�����;�!�9�d�f�f�W���	����l��B1�A݊�g�i�u�1�;�)��������l��hZ�Gʭ�'�4�
�:�$��ށ�P���F��X�����g�
�g�i�w�)�(�������P�������1�!�%�d�d�;�(��&���F��D�����%�6�;�!�;�k�F���s���C9��h��@���%�u�h�&�3�1��������AN��D�����8�
�`�3��k�(��Y�ƹ�@��R
�����;�!�9�c�f�t�}���Y����U��Y�����h�_�u�u�w�}��������EU�������8�
�f�'�0�i�O���P���A�R��U���u�u�u�4��2��������9F�N��U���d�d�6�&��(�N���	�����h�����0�!�'�'�$�'�_�������\��1��*��
�g�y�g�~�W�W���	����9��hW�*��i�u�!�
�8�4�(�������]��Y��3؊�
� �c�b�'�t�\ϫ�
����WN��h�����#�g�g�|�]�}�W���Y����l��C1��*��`�%�u�h�$�9��������G	��E�����<�;�1�%�$����@ù��J��G����u�:�d�3��i�G���Y����G��X	��*���!�'� �&�0�8�_�������R��E�����;�1�4�
�8�.�(���K���l�N��Uʥ�&�
�
�4�#�;�(��&���F��S1�����#�6�:�}�2�4�ǭ�����C	��h_�� ��b�%�|�f�~�f�}���Y����lW��B1�B���u�h�&�1�;�:��������F��P ��]���d�3�
�m��o�W�������V��G1�����9�d�
�|�l�}�W���YӖ��9��D�� ��e�
�d�i�w�)�(�������P�������&�2�0�}�8�o����M�ߓ�O�G����u�%�&�
�"�l�Nց�K���@��[�����6�:�}�;�>�3�ǘ�&���� ^��N�� ���2�0�}�%�4�3����H����]ǻN�����3�
�l�
�d�a�W���Y�����R	��*���c�f�%�u�?�3�_���&�ד�F9��1��]���h�r�r�u�;�8�}���Y���G��\�����m�
�f�_�w�}����
����9��h_�C���u�h�}�
�����Nù���������f�f�%�|�]�}�W�������]9��Q��M���%�u�h�}���F���&����l��V �����
�0�
�l�g�f�W�������@��h[�� ��c�
�g�i�w�/����&���� S��G\�����7�!�3�
�d�o����s���B��D�����3�
�e�m�'�}�J���&����l ��^�*��4�1�$�<������H���9F������2�
�
� �d�l�(��E����l��1��*��g�%�u�;�w�?��������^��d��Uʤ�
� �d�d��n�K���Y���F��D ��*���
�m�b�"�2�}����H����lW��1��]���h�r�r�u�;�8�}���Y���G��W�� ��e�
�f�_�w�}��������T��N�U���4�g�g�
�"�o�Nׁ�K����\��XN�N���u�'�d�3��k�(��E����^��1��*��
�g�4�1�#�-�B؁�����l��d��Uʧ�g�3�
�f�c�-�W��[����[����*��
� �g�f��l�JϿ�&����G9��1�U���0�w�w�_�w�}�(܁�����9��R��W���"�0�u�!�'�l�G�������
F�V�����
�#�d�e�w�1����[���F��1��*��b�%�u�h�u�� ���Yے��lW��h��*��c�h�4�
�8�.�(���H���V
��L�N���u�'��d�1��G���	�����h�����0�!�'�&�>�)����ۓ��Z��SF��*���&�
�#�a�d��1���?����uO��X1�����'� �&�2�2�u�G���Y����P��B1�Fӊ�d�f�x�u�8�3���P���9F���*ފ� �g�f�
�e�a�W���&����P9��T��]���;�1�!�%�o����Kʹ��F�D�����8�
�`�3��e�D���P��ƹF��h8��*���g�`�
�g�k�}��������E��X�����1�!�%�m��(�E��&���F��P ��]���
�b�3�
�o�j����B�����h��D��
�g�i�u�#�����&����\��_��*���=�}�;�<�9�9��������_��h]��3�������{�2��������]��Y��R��s�!�%�f��(�F��&���K��S�����|�|�|�_�w�}�(���H����CT�
N�����c�3�
�f�g�-�W���Y����_��B1�A܊�g�n�u�u�%�4�ށ����� 9��R��]���
�f�
� �f�m�(���ƾ�9��P1�E���_�u�u�
��o����J�Г�F�F����a�3�
�f�o�-�W����ԓ�F9��Z��G��u�u�'�<�>����J����Z���*���
�0�
�d�n�2�W���&����T��G\����u�
�
�a�1��E���	���N��G1�L���2�a�l�u�%�/�C���&����l��d��Uʧ�<�<�3�
�d�m����D�θ�C9��h��D��
�d�:�u��(�F��&���9F���D���
�`�e�%�w�`�_���&����U��X�����:�u�%�6�9�)����H��ƹF��R�����m�
�g�i�w�)���L����
Q��G]�����%�6�;�!�;�l�F��Y����V��Q��E���%�u�h�}�:��D؁����� 9����U���6�;�!�9�f�l�L���YӔ��9��h\�B���u�h�}�:�;�%�2�������R��h!��0���9�&�3�
�b�j�����ƭ�l��D��ۊ�|�_�u�u�2�e����O�ޓ�F�F����g�'�2�f�g�}����	����@��A_��\�ߊu�u�0�l�1��A���	���N��G1�A���
�c�l�%�w�2�W�������l
��h_����u�0�
� �f�n�(��E����^��Y�� ��g�
�f�-�%�<�(���
����9��d��Uʦ�9�!�%�e�1��C���	���l�N��Uʥ��9�
�
�"�l�Oف�Kӑ��]F��R�����3�
�a�l�'�u�^��^���V
��d��U���u�&�9�!�'����Iù��l�N�����%�d�3�
�c�n����D�θ�C9��h��D���
�f�-�'�6�����&����O��N�����!�%�g�3��i�N���Y���@��C��*���d�d�
�g�6�9��������l ��Z�*��n�u�u�&�;�)���&����A��h��G���
�g�i�u�#�-�Dց�����Q��EN�����'�2�f�g�~�W�W�������CW��Q��A���%�u�h�_�w�}�W���&����lU��B1�M܊�g�"�0�u�$�1����K����R��h�E���u�d�|�0�$�}�W���Y����V
��Z�*���d�g�
�f�]�}�W���&����9��h_�F���u�h�w�w� �8�Wǭ�����uT��R	��M��u�u�<�;�3�<�(���
����T��G�����u�e�n�u�w�.����	����W��E	��*���g�g�
�g�k�}����J����S��h����0�b�3�
�b�j����s���@��C��@Ҋ�0�:�2�;�1��A���	���N��[1�����
�0�:�2�9�;�(��J����\��Z��E���
�`�f�%�~�W�W�������CW��Q��A���%�u�h�}�2����&����S��G\�����8�
�
� �f�i�(��B�����h��D܊� �d�b�
�e�a�WǪ�	����l ��[�*��:�u�8�
�g�3����&����l��d��Uʦ�9�!�%�b�1��A���	���N��G1�*���d�a�
�g�6�9��������l ��X�*��n�u�u�&�;�)��������R��N�U���u�u�u��9�8�(���&����lW��B1�@܊�g�"�0�u�$�1����N����P��h�E���u�d�|�0�$�}�W���Y����V��B1�Fڊ�g�_�u�u�2����&����V��G]��H�ߊu�u�u�u�6�:�F�������\��B1�F܊�g�"�0�u�$�1����N����P��h�E���u�d�|�0�$�}�W���Y����l_��^1��*��e�%�n�u�w�.����	¹��lU��1��U��_�u�u�u�w��;���&����	��h�����
�c�l�%�w�5��������C9��h]�E���}�|�h�r�p�}����s���F�G1��%���:�
��9��2�(���	����F9��]��F�ߊu�u�0�
�:�o�(���K����CT�
N�����f�'�2�f�`�}����	����@��A_��\�ߊu�u�0�
�:�o�(���K����CT�
N�����3�
�e�f�'�}����
����A��V�\�ߊu�u�0�
�:�o�(���K����CT�
N�����f�'�2�f�`�}����
����A��V�\�ߊu�u�0�
�:�o�N�������]9��h]�D���u�h�}�8��m�(���J����CT��EN����d�3�
�a�c�-�^�ԜY�ƿ�_9��G\�����d�d�%�u�j�W�W���Y�Ƽ�e��h[�� ��c�
�f�"�2�}����J����lT��1��]���h�r�r�u�;�8�}���Y���C9��[\��*���
�l�f�_�w�}��������l��X�����
�a�l�%�w�`�_���&���� _��R�����3�
�a�d�'�}�Ϫ�	����l ��Z�*��n�u�u�&�;�)��������
T��N�U���u�u�u�&�;�)��������W��N�����&�9�!�%�n�9��������lT��1��]���h�r�r�u�;�8�}���Y���C9��[\��*���
�l�f�_�w�}��������U��W�����h�}�8�
��8�(��KӞ����T�����d�d�n�u�w�.����	�Г�F9��^��G��u�!�%�
�"�o�Gہ�KӇ����G1����c�|�_�u�w�8�(���KĹ��l^��h�I���u�u�u�u�#�-�F�������
9�������8�
�g�3��o�(��I���W����ߊu�u�u�u�'�>��������]ǻN�����8�g�
� �o�n����D�θ�C9��h��B���%�u�:�u�'�>�����ד�]ǻN�����8�g�
� �o�d����D�Ν�r(��y-��*���c�f�%�u�9�}��������U��]��G��u�u�&�9�#�-�(���J����CT�
N�����e�
� �f�c��EϦ�Ӈ��P	��C1��D��n�u�u�&�;�)��������W��N�U¦�9�!�%�l�%�:�D��Y����G��\�����m�d�%�|�]�}�W���&����9��C1��*��a�%�u�h��8�(���L����R��h����4�
�:�&��+�(���s���@��C��D���
�m�c�%�w�`�}���Y���C9��[\��*���d�g�
�g� �8�Wǭ����� V��B1�Aۊ�g�e�u�u�f�t����Y���F���*���g�
�0�
�n�m�}���Y����G��1��*��f�%�u�h��0�(��&����V��G]�����%�6�;�!�;�l�F��Y����V
��Z�*���d�`�
�g�k�}��������l��h]�@ʴ�1�&�9�!�'�o����A�Փ�O��N�����!�%�a�3��e�C���Y���F�N�����9�
�
� �f�o�(��������h��Fي� �d�`�
�e�m�W���H����_��=N��U���u�0�
�8�d����MŹ��l�N�����%�`�3�
�f��E��Yۏ��CW��B1�@���u�;�u�8��h����Jʹ��]ǻN�����8�f�
� �f�o�(��E����^��[�� ��f�%�u�'�#�-�Aׁ�����lW�� 1��\�ߊu�u�0�
�:�n�(���H����CT�
N�����l�3�
�e�n�-�W���Y����G��1��*��f�%�|�_�w�}��������U��]�����h�_�u�u�w�}����H����l	��D1�����e�b�%�u�?�3�_���&����9��h_�L���}�|�h�r�p�}����s���F�E��*���l�d�%�n�w�}��������l ��_�*��i�u�u�u�w�}�%���¹��_9��E��G���
�e�b�%�w�5��������CU��Q��D���%�}�|�h�p�z�W������F�N��Lߊ�d�3�
�d�f�-�L���Yӕ��l��1��*��l�%�u�h��8�O�������F��SN�����%�
� �f�g��E��Y����V
��Z�*���d�c�
�g�k�}����O¹��T9��Z�����%�6�;�!�;�l�F��Y����V
��Z�*���d�b�
�g�k�}����&����
Q��G\�����&�0�
�
�2��O��B�����h��A؊� �d�m�
�e�a�WǪ�	����A��W�U���u�&�0�
��8�(��@��ƹF��R����
� �g�a��n�K���Y���F��h8��G���3�
�g�a�'�}����Q����W��B1�Aۊ�g�e�u�u�f�t����Y���F������d�
�0�
�n�d�}���Y����G��1��*��c�%�u�h�]�}�W���Y����G��1��*��`�%�u�=�9�u��������l��X�����
�g�g�%��t�J���^�Ʃ�@�N��U���%��9�
�n�/���@��ƹF��R����
� �g�c��o�K�������
9��P1�B���:�u�%�6�9�)����H��ƹF��R����
� �g�b��o�K�������l ��\�*��4�1�<�8�e�/���K����F�D�����b�3�
�c�f�-�W��Q���� 9��h\�D���u�:�u�%�4�3����H���9F���*���a�
� �g�f��E��Y۔��9��h\�B���u�;�u�0��0�C؁�����9��UךU���0�
�8�a��(�E��&���F��X������!��0�#�/�8�������@9��h\�B���u�;�u�6�'�j��������_��G�U���&�9�!�%��(�D��&���FǻN��U���
�
�0�<�3�4�(���Y����N��[1��ي� �f�e�
�e�m�W���H����_��=N��U���u�0�
�8�f�;�(��L����9F���*���`�
� �g�c��E��Yے��l^��Q��@���%�u�;�u�2����&����U��G\����u�0�
�8�b����L����Z���*���d�m�1�8�%�<�(���K����CT��X�����;�!�9�d�f�f�W���
����^��h��G��
�g�i�u�#�-�Oށ�����^��Y
�����8�`�
�0��l�E��Y����V
��Z�*���g�l�
�f�k�}�W���Y����C9��Y�����g�"�0�u�$�1����A����lR��F�U���d�|�0�&�w�}�W���YӇ��P	��C1��F���_�u�u�0��0�Bہ�����9��R�����u�u�u�0��0�B܁�����9�������'�6�;�d�1��@���	����[�I�����u�u�u�u�w�-����&����l��=N��U���
�8�`�
�"�o�F܁�J���9F�N��U���6�;�!�9�d�n� ���Yە��l��\�� ��m�
�g�e�w�}�F�������9F�N��U���6�;�!�9�d�k�}���Y����G��1��*��l�%�u�h��0�(��&����W��G\�����%�6�;�!�;�l�F��Y����V
��Z�*���f�a�
�g�k�}����H�ד�F9��Z��Gʴ�1�&�9�!�'�k����M�ߓ�O��N�����!�%�m�3��i�@���Y���@��C��Fӊ�0�:�2�;�1��C���	�ƴ�AF��h�����#�
�|�_�w�}��������U��X�����h�}�8�
�g����Kʹ������*���`�
� �f�b��E��Y����V
��Z�����a�l�%�u�j�u�����ߓ�F9��Z��Gʴ�1�!�%�c��(�F��&���9F���*���c�
� �f�`��E��Yە��l��Z�����'�4�
� �d�k�(������C9��Y�����d�n�u�u�$�1����H���� R��h�I���!�%�d�f�1��C���	�ƭ�WF��[1�����3�
�a�`�'�t�}���Y����G��1�����4�
� �g�o��E��Yے��l��R	��M��:�u�6�%�%�:�D��P���F��[1��܊� �f�g�
�e�a�WǪ�	����l��h]�Dʴ�1�'�#�
�"�n�B؁�K��ƹF��R�����3�
�a�e�'�}�J�ԜY���F��G1�*���d�f�
�d� �8�WǪ�	�ӓ�F9��X��G��u�u�d�|�2�.�W���Y�����T�����g�
�n�u�w�.����	˹��lW��1��U��}�8�
�
�"�l�Eف�KӞ����T�����d�d�n�u�w�.����	�Г�\��B1�Eӊ�g�i�u�&�;�)��������W��N��ʴ�
�:�&�
�!��^�ԜY�ƿ�_9��GW�� ��d�
�g�i�w��6���7����T9��\�����0�
�8�m�1��C���	����F�D�����3�
�c�e�'�}�J�������9��h]�A���u�;�u�0�o�/���M����F�N�����8�
�
�4�#�;�(��&���F��S1�����#�6�:�}�2�4�ǭ�����@��Z��*���b�d�%�|�d�t�L�ԜY�ƿ�l��h_�� ��d�%�u�h�]�}�W���Y����V��B1�L���u�=�;�}���>���H����_��G\��\��r�r�u�9�2�W�W���Y�Ƹ�C9��h��B���%�n�u�u�w�}��������@��B1�G؊�d�i�u�!��2����������^�����0�}�=�4�#�;�(��L����U��UװU���&�
�8�
�"�l�Fځ�J���9F�N��U���
�
� �d�g��Eϩ�����f'��~ �����f�`�}�|�j�z�P������F�N�����f�3�
�g�g�-�L���Yӕ��]9��D��*ۊ� �d�m�
�d�a�W���Y�����hY�����l�a�%�u�?�3�_���&����9��h_�G���}�|�h�r�p�}����s���F�D�����d�3�
�l�`�-�L���Yӕ��]9��D��*ۊ�:�
� �g�c��E��Yە��]9��D��*ۊ� �d�m�
�d�%�Ͽ�&����G9��1�N���u�&�2�
�$�4����&����l��S��U���u�u�!�%�d����L˹����YN�����8�g�
� �e�e�(��I���W����ߊu�u�u�u�2����&����Q��G\�U���&�2�
�&�>�3��������R��N�U¦�2�
�&�<�9�;�(��N����K	��V�����
�#�
�|�]�}�W�������U��^�����h�%��9��j����K�ޓ�N��
�����f�|�_�u�w�0�F߁�����9��R��]���'�9�"�d�1��G���	�ƣ���Y1�����
�
�:�
�"�o�C߁�K��ƹF��Z�*���g�c�
�g�k�}��������A��^�U���u�0�
�8�c����O����]ǻN����
� �g�m��o�K�������T��C1�����a�`�u�'�#�-�@؁�����9��UךU���8�d�
� �d�h�(��E����^��1�����4�
� �f�c��EϦ�Ӈ��P	��C1��D��n�u�u�!�'�i����H�ד�F�F�����0�e�1�8�%�<�(�������T��N��U���
�a�3�
�f�l����s���G��1��*��f�%�u�h��0�E�������T��Q��F���%�u�:�u�'�>�����ד�]ǻN����
� �f�`��o�K�������T��h
�����;�<�
� �d�o�(���Ƹ�C9��h��F��
�g�n�u�w�)��������P��N�U���
�:�<�
�2�)�ǫ�
����WN��a��*���'�2�a�g�~�v��������C9��g�����;�&�2�|�]�}�W���H����S��h�I���9�
� �d�c��FϿ�Ӕ��l ��[�*��n�u�u�!�'�e�(�������G9��h[�*��i�u�u�u�w�}��������_��h\�����}� ����;�(��&���F�_��U���0�_�u�u�w�}��������EW��UךU���8�g�b�1�:�/��������9��R��]���
�f�
� �f�n�(���ƿ�_9��G]�����f�g�|�_�w�}���A����G9��D�� ��b�%�u�h�]�}�W���Y����\��h��G��"�0�u����9���&����
U��F�U���d�|�0�&�w�}�W���YӇ��P	��C1��D؊�n�u�u�!�'�d�(�������l ��Z�*��i�u�%�f�����M����	��U�����e�1�8�'�6��(���K����CT�=N��U���g�c�1�8�%�<�(���J����CT�
N��*���<�
� �f�f��Eϱ�Y����A��1�����4�
�d�3��l�E���P���F��G\�*���:�2�;�3��n�@���Y���C9��h�����g�g�%�u�%�?�����֓�V��P��؊� �f�g�
�e�f�W�������U�� ]�����h�}�0�
�:�l�(���H����CT��EN�����%�e�;�!�1��@���	����F�C��*���g�b�
�g�k�}��������G9��P1�B���;�u�0�
�:�o�(���K����CT�=N��U���a�3�
�d�g�-�W��Q����U
��h��G��
�g�:�u�>�3��������G9��h\�A���|�_�u�u�:�h����K�ғ�F�F�����0�3�
�d�a�-�W���Y����G��1��*��l�%�|�_�w�}��������U��N�U¡�%�m�
�0�8�:����&����l��O�����:�&�
�#��t�}���Y����l ��^�*��i�u�9�
��(�N���	�ƭ�WF��A\�� ��d�%�|�_�w�}��������S��N�U¦�9�!�%�`�%�:�D��Y����V
��Z�*���
� �d�e��o�L���YӒ��
9��h_�D���u�h�}�0�$�:����H����^��h����&�9�!�%�g�;�(��I����l�N����e�3�
�a�n�-�W��[����[�������4�0��'�4�(���A����lR��N�����:�&�
�#��t����Y���9F���*��
� �f�g��o�K���H�ƻ�V�B,�����&�
�!� �#�/�(��&����W��S�����;�!�9�f�e�}����[����F�C��D���3�
�a�l�'�}�J���[ӑ��]F��u1��*���0��'�6�"�8�F�������W��
N��*���&�
�#�
�~�8����I��ƹF��Z��Eي� �f�f�
�e�a�W��Y����N��h��6���
�!� �!�%��Cׁ�����R������!�9�f�c�w�1����[���F��G1�@���
�c�`�%�w�`��������l��C�����/�}�;�<�9�9��������l*��G1�����a�l�y�a�~�W�W�������9��h]�A���u�h�w�w� �8�Wǭ�����Q��1�Aӊ�e�u�u�<�9�9����)����W9��h��\���9�0�w�w�]�}�W���&����U��\�����h�%�&�
�"�l�N߁�K����W	��C��D��u�u�!�%�f�e����N�ߓ�F������,� �
�e��(�D��&���F��@ ��U���_�u�u�8��m����K�ד�F���*���<�
�0�!�%�.����������Y������3�
�d�o�-�^ê�&����T��B �����}�e�u�u�:��(���H����CW�C����!�u�|�|�~�W�W�������9��h_�G���u�h�%�&��(�F��&���F��@ ��U��n�u�u�!�'�l�B���&����l��S�����3�
�a�e�'�u�FϺ�����W�=N��U���
�d�
� �a�d����Dӏ��T9��1��*��
�d�c�u�w�}�������9F���*��
� �c�d�'�}�JϷ�����9��hX�*��`�u�u�u�8�3���B�����h_�*���b�l�%�u�j�0����O����Q��G]��M���d�1�"�!�w�t�}���Y���G��_�� ��c�
�d�i�w�)�(�������P�������&�2�0�}�:��G���&����l��]�\�ߠu�u�!�%�f�m����Lƹ��Z�C��A݊� �b�l�%��e�Z������\F��d��Uʡ�%�d�d�3��k�(��E�Ƹ�C9��h��B���%�}�m�x�f�9� ���Y����F�C��D���3�
�m�
�d�a�W���&����U�� ]��F¡�
�;�0�0��3����ے��lP��T��*���b�`�%�|�w�2��������G��EF�����0�}�8�
�`�>��������l��G�����}�:�<�!�0�/��������G��Y�����3�
�m�
�f�t�J������\9��C�� �&�2�0�}�:��@���
����lQ��h�\��f�u�9�0�u��}���Y����T��Q��Gي�d�i�u�8��h����H¹��P�_�����:�e�n�u�w�)���M����U��G]��H�ߊu�u�u�u�'�>�����Г�F��R �����`�
� �m�`�-�_���D����F��D��U���u�u�%�:�f�;�(��&����F�C��D���3�
�a�
�f�a�W���&����P9��T��]���<�0� �&�0�8�_���&����U��]��F���a�|�_�u�w�0�(��&����S��N�U���
�:�<�
�2�)�ǭ�����V ��B �����}�%�6�;�#�1�Bہ�?����u ��q(��\ơ�
�;�0�0��3��������@��Z��Gߊ� �m�d�%��l�FϺ�����O�G�U���!�%�d�b�1��Bށ�K�����h_�*���m�`�%�u�8�}��������ES��(��3������|�]�}�W���&����U��^�����h�%��9�����@ƹ��W��S�����b�n�u�u�#�-�F݁�����9��R�����9�2�6�#�4�2�_�������U��Y�����!�%�d�
�"�l�Aׁ�H�ʸ�l��R	��]���<�;�1�r�p�{��������@��B1�G؊�d�f�x�u�8�3���P���9F���*��
� �d�e��l�K���&����l_��B1�Lߊ�f�d�x�d�3�*����P���F��G1�D���
�m�f�%�w�`��������U��\�����b�1�"�!�w�j�L���YӒ��lW��h��M���%�u�h������N����W��X����n�u�u�!�'�l�D���&����CR�
N����
� �l�`�'�u�FϺ�����O��N�����d�`�3�
�`��D��Y����lW��B1�B���}�d�1�"�#�}�F��Y����^��Y�� ��d�
�f�i�w�2�E�������9��_����!�u�d�n�w�}����H�ޓ�F9��Y��F��u�:�d�d�1��C؁�K����W	��C��D��u�u�!�%�f����@ù��Z�_�����u�&�2�0��0�(݁�����9��N����0�}�%�6�9�)���&�����RN��W�ߊu�u�8�
�c����Jù��Z�G1��؊�b�3�
�g�o�-�_���Y�ƨ�D��^����u�8�
�a��(�E��&���F��a��*���3�
�g�m�'�u�DϺ����� U�=N��U���
�a�
� �e�i�(��E�Ƽ�e��h\�����g�m�%�}�g�9� ���Y���9F���*��
� �g�d��n�K���&����lR��Q��@���%�}�f�1� �)�W��B�����h_�*���g�b�
�f�k�}����&����|��p������
�$�4�����LĹ��@��X������!��0�#�/�8�������9��h\�@���|�_�u�u�:��C���&����CW�
N�����
� �a�b�'�u�E��Hӂ��]��G�U���!�%�d�e�1��N���	��� ��h��9��� �
� �!�'�$�F���/����^��h�G���u�u�:�;�8�m�L���YӒ��lW��h��G��
�d�i�u�/��:��� ����~��^��*��
�
� �g�`��E��Y����W	��C��\�ߊu�u�8�
�b�;�(��O����[��C
�����
�0�!�'�"�.����Q�ԓ�V��Z�U���;�<�;�1�6�����&����l ��G�U���!�%�d�f�1��A���	�����h^��G���$�}�d�x�f�9� ���Y����F�C��D���3�
�c�l�'�}�Jϼ��֓�R��F^��Dʱ�"�!�u�d�l�}�WϪ�	����l ��X�*��i�u� �
��o�N���Q����\��XN�\�ߊu�u�8�
�a�;�(��I����[�L�����}�<�;�1������A���F��P ��]���6�;�!�9�f��@�������V�=N��U���
�b�3�
�b��E��Y����_	��T1�����}�;�<�;�3��(���L�Փ�O������1�4�
�:�$�����?���l�N����
� �`�d�'�}�J���[ӑ��]F��^	��¡�%�d�
� �b�h����Gӕ��]��V�����
�#�g�f�~�}����[����F�N�����d�
�4�!�1��D���	�����h�����0�!�'�'�$�'�_�������^��1��*��c�%�|�f�~�f�}���Y����_��B1�A܊�g�i�u�e�w�5����&����_��h��D��
�g�h�4��2�����ғ�F��D��D��u�u�!�%�f�;�(��H����[�L�����}�;�<�;�3�.�(���&����W��G]��Iʠ�&�2�0�}�'�>��������^������w�_�u�u�:��G���&����l��S�����
� �d�l��n�E���Y�ƨ�D��^����u�8�
�d�1��D���	�����h�����0�!�'�'�$�'�_���������V�����
� �d�b��o�[��P���F��G1�*���`�f�%�u�j�.��������V��EF�����0�}�8�g�f�>��������F9��1��\��� �&�2�0��%�(�������l��UךU���8�
�f�3��h�A���Y���D��_��]���;�1�%�&��(�F��&���F��P ��]���6�;�!�9�f��A�������V�=N��U���
�a�3�
�e�j����DӒ��lW��Q��G���%�}�a�x�f�9� ���Y����F�C��Gߊ� �d�f�
�f�a�W���&����P9��T��]���<�0� �&�0�8�_���H����G9��h_�@���|�`�|�n�w�}����KŹ��lW��1��U��!�%�d�
�"�l�@݁�K����F��S�����|�_�u�u�:��@���&����l��S�����:�<�
�0�#�/��������[��^	��¸�;��3�
�f�e��������G��EF�����0�}�e�u�w�0�(������� P��F�X���:�;�:�e�~�t�L���YӒ��lT��Q��@���%�u�h�w�u�*����
����WN��D\�� ��l�
�g�u�w�4��������]��[�*��|�0�&�u�g�f�W�������
9��h_�@���u�h�8�;��;�(��A����G	��Y�����;�<�;�1�#�-�Fց�����F9��_��D���1�"�!�u�8�4����ۓ��Z��SF����
�4�!�3��n�F���P����[�������2�'� �&�0�8�_���&�ߓ�R��Q��F���%�|�k�u�w�3�W�������V��Y�����!�%�d�
�6�)����J�ד�O�
[�U���0�w�w�_�w�}����&����V��G\��Hʦ�1�9�2�6�!�>��������V��1����a�|�~� �$�:����	����@��A_��3���|�_�u�u�:��G���&����l��S�����:�<�
�0�#�/�����ι�@��R
�����6�&�
� �f�m�(��U���l�N����
�:�
� �f�k�(��E����^��1��*���c�%�u�:�w�-��������lW�=N��U���
�d�3�
�a�m����D������YN�����g��d�3��h�E���Y�ƭ�l��D�����e�u�9�0�u��}���Y���� T��B1�AҊ�g�i�u�d�w�5�����ԓ�F9��W��G��4�
�:�&��+�E��PӃ��VF�UךU���8�
�f�3��l�A���Y���G��D1����f�u�'� �3�/�������� T��G�U���!�%�f�
�"�o�Bׁ�K���4��P�����:�0�
�
��h����J����K	��V�����
�#�
�|�]�}�W���&�ӓ�F9�� 1��U��!�%�d�
�"�h�B���Q���F��@ ��U���_�u�u�8��k����H�֓�F�F�����'�2�f�d�w�2�W�������l
��h_����u�8�
�b�1��Cށ�H���@��[�����6�:�}�0�>�8��������V��C��#���3�
�f�
�c�q�E���s���G��V�� ��`�%�u�h��-��������lW���*��
� �c�d�'�t�}���Y���� _��B1�D���u�h�w�w� �8�WǪ�	����l ��_�����u�%�6�;�#�1�A܁�PӃ��VF�UךU���8�
�
� �f�l�(��E�ƿ�W9��P�����:�}�;�<�9�9��������_��h_�U���;�<�;�1������A���l�N����
� �c�l�'�}�Jϭ�����Z��R�� �&�2�0�}�e�l����AĹ��F�B �����}�%�6�;�#�1�F݁�?���9F���*���3�
�e�
�e�a�W���&����P9��T��]���<�;�1�4��2�����ԓ�O������1��
�
�"�k�@���P��ƹF��Z��G���
�g�
�g�k�}�F������uT��h��C���%�u�u�%�4�3����H����F��D��E��u�u�!�%�c����J����[�L�����}�;�<�;�3�.�(���&¹��lQ��h�U���;�<�;�1�6�����&����lU��N�����e�n�u�u�#�-�Cہ�����l��S��U���u�u�4�
�8�.�(���&����[����*���3�
�c�
�e�m�W���H����_��=N��U���u�
�%�3��j�(��s���G��[�� ��l�%�u�h�u�� ���Yۓ��Z��SF��*���
�
� �b�f�-�^������]��V�����
�#�g�d�~�}����[����F�C��A܊� �b�`�%�w�`��������l��C�����/�}�;�<�9�9��������P��h��B���%�|�`�|�l�}�WϪ�	����U��W��G��u�!�
�:�>�����ە��U��^	��]���;�1�8�;��k����N����J��h�����}�;�<�;�3�z�P�������9��hY�*��f�x�u�:�9�2�G���P��ƹF�N�����m�3�
�`��l�K�������T��A�����0�<�0�&�0�8�_���&����U��W��D���g�|�_�u�w�)���&���� T��G_��Hʦ�1�9�2�6�!�>����������^	��¡�%�a�
�0��e�O��M����F�C��A���
�d�d�%�w�`�_�������l
��h_��U���
�a�'�2�d�o�^�ԜY�Ƹ�C9��h��B���%�u�h�&�3�1��������AN��^�����}�;�<�;�3�)���&����_��G�����!�2�'� �$�:����I���@��Z��*���!�3�
�d��l�D��Y����G	�G��\�ߊu�u�8�
�f�;�(��&���F�N�����&�2�0�}�:��G���&����CT�	N�����}�%�6�;�#�1�F݁�O����_��^�����u�8�
�g�1��D���	�����h�����0�!�'�&�>�)����Q����T�������!�9�`�
���1���?����J��h�����}�;�<�;�3�z�P�������
9��h_�@���}�d�d�1� �)�W���P����F�C��@ي� �b�l�%�w�`��������l��C�� ���2�0�}�g�f�;�(��&���F��D�����%�6�;�!�;�l�(���P��ƹF��Z��A���
�e�
�g�k�}�F������@��R
��G���3�
�m�
�e�}�W�������C9��Y����
�d�|�0�$�}�G��Y����^��1��*��
�g�i�u�#�����&����\��Y������
�
� �a�j����Rӓ��Z��SF��*���&�
�#�g���^�ԜY�Ƹ�C9��h��M���%�u�h�w�u�*����
����WN��G1�*���m�d�%�|�i�.����Q����\��h��G��|�u�9�0�u��}���Y����Q��B1�F���u�h�w�w� �8�WǮ�+����G9��Q��@݊�g�h�4�
�8�.�(���M���V
��L�N���u�!�%�`��(�F��&���F��Z��G���
�f�m�%�w�2�W�������l
��1��3�������~�W�W�������l ��V�*��i�u�!�
�8�4�(�������V��RF�����0�}�7�4�$�:�(܁�����9��B�\��u�u�!�%�b�;�(��O����[�L�����}�g�'�2�d�i�W���	����@��A_��D���0�&�u�e�l�}�WϪ�	����U��[��G��u�!�
�:�>�����ۓ��Z��SF����
�4�!�6�$����N����M��Y�����0�%��d�1��Cځ�K����F�C��Cۊ� �l�b�%�w�`�U���������Y�����
�
� �l�`�-�^��
����WN��h�����#�g�f�|�w�1����[���F��G1�*���l�b�%�u�j�.��������V��EF�����}�;�<�;�3�-�ށ�&����l ��[�����`�|�n�u�w�)���&����
W��N�U���
�:�<�
�2�)�ǭ�����Z�������8�;��c�1��@܁�J�ʸ�l��R	��]���<�;�1�r�p�{����O����l_��h�F���u�:�;�:�g�t�^��Y����^��1��*��m�%�u�h�'��݁�&����^��G]��Fʱ�"�!�u�f�l�}�WϪ�	����U��\�����h�w�w�"�2�}�����μ�@T��h��L���%�|�i�&�0�8�_�������l
��1�\���9�0�w�w�]�}�W���&�Г�F9��W��D��u�!�
�:�>�����۔��Z��B �����}�:�g�d�4�.�(���@�Փ�O�G����u�u�u�8��j����&����S��N�U���
�:�<�
�2�)�Ǭ�
����@��R
�����f�3�
�b��o�[��P��ƹF��Z��B���
�f�c�%�w�`��������U��V�����u�u�u�:�9�2�G��Y����^��1��*��d�%�u�h�u�� ���Y۴��T��a1�����e�f�%�u�w�-��������9�������w�_�u�u�:��O�������W��h�I���!�%�c�
�"�l�E؁�KӞ����T�����d�d�n�u�w�)���&����_��G\��H���w�"�0�u�'�.�(ށ�����l��
N��*���&�
�#�g�d�t����Y���9F���*܊� �`�f�%�w�`��������l��C�����/�}�;�<�9�9��������l ��_�����d�|�n�u�w�)���&����
S��G\��H���4�2�d�4�;�2����&�ד�9��h_�L���u�:�u�%�4�3����H���9F���*���3�
�g�d�'�}�J�������l��h]�Bʺ�u�;�0�3�8��(���&����]ǻN�����g�3�
�e�f�-�W��Q����T9��E��F��u�:�u�%�4�3����H���9F���*���3�
�f�g�'�}�JϮ�/���� 9��h_�C���}�f�1�"�#�}�D��Y����^��1��*��d�%�u�h�u�� ���Yە��]��G1��؊�c�'�2�a�e�t�Iϭ�����R��X ��*���a�e�|�0�$�}�G��Y����^��1��*��m�%�u�h�$�9��������G	��E�����;�<�;�1�&������ӓ�F9��\��G���a�|�_�u�w�0�(�������P��N�U»�"�<�;�<�����N˹���������!�9�d�d�l�}�WϪ�	����U��]�����h�}�<�;�>�����I����\��G1�����9�d�d�n�w�}����N˹��lT��1��U��w�w�"�0�w�.����Q����_T��1��*���l�%�|�k�$�:����	����@��A\��E���0�&�u�e�l�}�WϪ�	����U��X�����h�}�7�:������&����G��x�����
�
� �g�b��E�������K!��x��2���!�'��
�&�<�(ށ�����9��N�����
��e� ��/����&����B��h�� ��d�
�g�n�w�}����N����V��G_��Hʼ�0�
�
� �c�j����J�����Y��E��u�u�!�%�o����@����Z�_�����u�!�%�b��(�E��&�����T�����f�`�u�9�2��U�ԜY�Ƹ�C9��h��G��
�g�i�u�f�}����Q����_��B1�Cي�a�h�4�
�8�.�(���&����_��^�����u�8�
�g�1��Nց�M���G��\�� ���f�%�}�d�3�*����P���F��G1�*���g�e�
�g�k�}�F������G�� W�� ��c�
�a�h�6�����&����O��[��W���_�u�u�u�w�0�(�������_��N�U���
�:�<�
�2�)�Ǭ�
����@��R
��*���g�m�3�
�`�m����K���9l�N��Uʡ�%�m�
� �e�n�(��E�ƿ�W9��P�����:�}�0�<�2�.����Q����_T��h��G���
�f�y�c�~�W�W���Y����^��1��*��f�%�u�h�$�9��������G	��E�����<�;�1�%��1�(ځ�N����Q��h�Y��|�_�u�u�w�}����AĹ��lT�� 1��U��&�1�9�2�4�+����Q����I��^	��¥��9�
�m�1��@���	���O�=d��U���u�!�%�m��(�E��&���F��S1�����#�6�:�}�2�4�ǭ�����C9��g�����;�&�2�y�`�t�}���YӒ��l^��B1�Fߊ�g�i�u�d�w�5��������V��_1�����
�g�`�%�~�a��������R��X ��*���g�f�|�u�;�8�U���s���G��_�� ��a�
�d�i�w�)�(�������P������� �&�2�0��?��������U��]�����f�|�n�u�w�)���&����P��G\��H���0�&�2�7�#�n����I�ԓ� F��EN��*���&�
�#�
�~�W�W�������l ��^�*��i�u�!�%�f�i����M����K	��V�����
�#�
�|�]�}�W���&�ғ�F9��_��G��u�&�2�7�#�l����M����K	��V�����
�#�
�|�]�}�W���&�ӓ�F9��\��D��u�!�
�:�>�����۔��Z��B �����}�7�4�&�0��(���J����CT�\��N���u�!�%�l��(�D��&���F��R�����!�a�3�
�e�l�����ƭ�l��D��ۊ�|�_�u�u�:��@���&����l��S�����d�d�'�2�c�m�W���Y����\��h��*���_�u�u�8��e����J�֓�F�F�����!�g�'�2�c�j�W���Y����\��h��*���_�u�u�8��d����J�ӓ�F������
�0�8�d�g�;�(��I���� W��X����n�u�u�!�'�d����K�ѓ�F���*���<�
�0�!�%�/����Q����T�������6�&�
� �f�o�(��U���l�N�����8�'�4�
�"�l�@݁�K�����hY�����f�g�%�u�%�.����	�ӓ�F9��V��G��u�u�!�%�1��C���	���N��G1�����4�
� �d�`��EϦ�Ӈ��P	��C1��D��n�u�u�!�'�.����JĹ��Z�_�����u�!�%�b�1��Gށ�H����C9��Y����
�|�0�&�w�m�L���Yӓ��P��V��&���6� �0�d�o�>��������9��R�����9�2�6�#�4�2�_�������]��Y�� ���&��&�
�#�(����&����A��_�\��|�_�u�u��>�(�������F��E��AҊ� �g�g�
�d�a�W���Y�����h��@ߊ� �g�d�
�d�*��������]��B1�MҊ�g�e�u�u�f�t����Y���F���*���`�
� �g�g��D�ԜY�ƹ�G9��h\�D���u�h�w�w� �8�Wǫ�
����WN��G1��&���!��&�9�#�����&�ѓ�l ��Z�*��u�u�;�<�9�9����8����F��U�� ����9�0�l�����M����O��[��W���_�u�u�;�2�;����&����U��G\��H���<�;�4�&�0��(���H����CU��Y
�����2�l�
�d�1��G���	����F�B �����"�g�3�
�c�n����D�θ�CT��h
�����;�3�
�a�`�-�W���Y����Q��E��A��|�_�u�u�9�8����&����G9��h\�L���u�h�}�8�f����Aǹ��	��G1�*��� �g�a�
�e�f�W�������U
��h]�� ��c�
�g�i�w�.�����ד�V��\����!�%�f�3��l�C���P���F��S�����f�;�!�3��l�@���Y���G��1��*��d�%�u�'�'�n�(�������U��G�U��� �1�'�9� �i����J�ߓ�F�F�����!�g�'�2�c�j�W���Y����9��h]�F���|�_�u�u�9�8����&ǹ��G9��h]�C���u�h�}�8�f����Lù��	��G1�*���3�
�g�g�'�t�}���Y����A ��@1��*��g�%�u�h��4����
����U��V�����;�u�'�0�0�d�(�������9��U�����0�4�n�