-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��LӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ��`�a�c��}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e�e�o��w�	�(���0����p2��F�U���;�:�e�n�w�}��������}F��s1��2���_�u�u�
����������}F��s1��2���_�u�u�
��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�Ƽ�9��V�����u������4�ԜY�Ƽ�F��~ ��!�����
����_������\F��d��Uʥ�d�4�
�9�w�}�9ύ�=����z%��N����o��u����>���<����N��
�����e�n�u�u�'�o��������z(��c*��:���n�u�u�%�c�m���Cө��5��h"��<������}�f�9� ���Y����F�G1��E���e�4�
�9�w�}�"���-����t/��=N��U���
�
�
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ғ�l��h�����o������0���s���C9��1��D��������4���:����U��S�����|�_�u�u���(���&����_�!��U���
���n�w�}����H����\��b:��!�����
����_������\F��d��Uʥ�a�d�0�d�6�����Y����`2��{!��6�ߊu�u�
�
�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����9��h��U���������}���Y����F��~ ��!�����
����_������\F��d��Uʥ�`�d�4�
�;�}�W���*����|!��d��Uʥ�c�e�0�e�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����9��1��*���u�u� �u���8���B�����h_��*���u� �u����>���<����N��
�����e�n�u�u�'�k�F���I����E
��N��!ʆ�����]�}�W���&ù��F��x;��&���������W��Y����G	�UךU���
�
�
�
��-����Cө��5��h"��<��u�u�%�c�f�8�F��6����g"��x)��*�����}�d�3�*����P���F��1�����4�
�9�u�w��W���&����p]ǻN��*Ҋ�
�
�u�u��}�#���6����e#��x<��F���:�;�:�e�l�}�WϮ�A�֓�lV��G1����������4�ԜY�Ƽ�9��R1�Oʚ�������!���6���F��@ ��U���_�u�u�
���(߁�	����\��b:��!�����n�u�w�-�O������)��=��*����
����u�FϺ�����O��N�����e�0�d�4��1�W���,�Ɵ�w9��p'�����u�
�
�
��}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y����l^��h��*���#�1�o����3���>���l��SUװ���=�!�6� �2�?�����ơ�u_��V��*���&�_�u�u�#�/����Y����l!��r<��<�����u�u���0�ԜY�ƭ�G��B��6���
������>���Y����V��T�����!�6� �0�>�W�W�������R��Q1����<�
�e�`�c�&�;���7����g?��
��Y���
�� �
���J���5����c3��q'��1��������%���Ĝ����V�DƝ�������<��W����V��{=��;���
���:�?�/�[���&����p*��|S�[��`�e�����;���J�ʄ�`9��y1��!׻�;�y��
���2��U����`?��s=��LƝ�����j�h�DÖ�*����l*��
V�C���_�u�u�:�$�<�Ͽ�&����G9��P��D�������g�W��B�����D��ʴ�
�:�&�
�8�4�(���Y����)��tN�U��n�u�u�6�9�)����	����@��Q��E��������4���Y����\��XN�U��w�e�w�_�w�}��������C9��h��*���
�u�u����>���<����N��S�����|�o�u�e�g�f�W�������R��V��!���f�3�8�g�m��3���>����v%��eN��U���;�:�e�u�j��G���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�l�F��*����|!��h8��!���}�u�:�;�8�m�W��[����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)����I����g"��x)��*�����}�u�8�3���Y���D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����W��d��Uʶ�;�!�;�u�'�>�����ԓ�\��c*��:���
�����}�������	[�^�����u�:�&�4�#�<�(���
����9��N��1��������}�FϺ�����O�
N��E��u�u�6�;�#�3�W�������l
��h_��U���
���
��	�%���Y����G	�N�U��w�_�u�u�$�:����	����U��N��1��������}�EϺ�����O�
N��E���_�u�u�!�%�?����
����P	��Y	��U���<�2�_�u�w�)�����ƪ�^9��T�����3�4�
��1�0�Mϭ�����Z�Y��W�ߊu�u�<�;�;�<�(���&����l5��D�����e�o�����4�ԜY�ƿ�T�������7�1�d�u�w��;���B�����Y�����e�<�
�<�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4����	�֓�l��A�����<�u�u����>��Y����Z��[N��E���4�
�9�
�%�:�Mύ�=����z%�
N��R�ߊu�u�<�;�;�-�G�������TF��d:��9�������w�n�W������]ǻN�����9�%�e�d�'�8�W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��P ��U���
�
�%�#�3�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�m�F���&����C��T��!�����u�h�p�z�}���Y����R
��h_�����2�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�H����TF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���&�2�4�u����������@��N��1�����_�u�w�4����	�ד�C9��S1�����u��
���}�J���^���F��P ��U���
�;�&�2�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������lT��E��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��n�u�u�&�0�<�W���&����_��Y1���������W�W���������h�����%�0�u�u���8���Y���A��N�����4�u�
�
��3����Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*ߊ�
�'�2�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�f�W���
����_F��1�����9�
�;�&�0�g�$���5����l�N�����u�
�
�
�'�+��������`2��{!��6��u�e�n�u�w�.����Y����9��h��U����
�����#���Q����\��XN�N���u�&�2�4�w��(ށ����5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���;�9�%�`�f�<�(���&����Z�=��*����n�u�u�$�:����&ƹ��R��[
�����o������M���I��ƹF��^	��ʴ�
�<�
�1��o�W���6����}]ǻN�����9�<�
�<��/�;���&˹��U��]��G��������4���Y����\��XN�N���u�&�2�4�w���������\��h_�����`�u�u����>���<����N��S�����|�_�u�u�>�3�Ͽ�&����P��h=�����3�8�d�o���;���:���F��P ��U���&�2�7�1�f�k�MϜ�6����l�N�����u�8�
� �d�d����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���
�c�u�u���8���&����|4�N�����u�|�_�u�w�4��������\��h��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϸ�&����\��X��Gي� �a�f�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����U5��C1�����:�
�f�'�0�h�N��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������:�
�:�%�e����I����	F��s1��2������u�d�}�������9F������3�
�!��%�����L����lS��T��!�����
����_������\F��d��Uʦ�2�4�u�
��(����H����lW��B1�D���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���
����@��d:��ي�&�
�u�u���8���B�����Y�����<�
�1�
�a�}�W���5����9F������2�%�3�e�1�l����Nʹ��l��RN�&������_�w�}����Ӗ��l��Q��D���e�g�3�
�c��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���3�'�d�0�f�l����Lƹ��\��c*��:���
�����l��������l�N�����u�
�
� �1�/�F���H�ԓ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w��(�������l��h_�� ��l�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Q��R��*���
�
� �a�a�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1�����0�
�
�
�����J����	F��s1��2������u�d�}�������9F������%�c�7�3�2��(���&����lR��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�e��������V9��1��*��
�f�o����0���/����aF�N�����u�|�_�u�w�4����	�ޓ�F ��E1�����g�3�
�e��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��hV�� ���'�d�0�d�f�;�(��&���5��h"��<������}�f�9� ���Y����F�D�����
�
� �3�%�l����K����W��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%��(߁�&¹��lU��h�����!�o�����4�ԜY�ƿ�T��	��*���
�
�
� �d�d�������5��h"��<��u�u�&�2�6�}����&ù��9��h]�*���'�4�,�o���;���:���F��P ��U���
�
�
�
��(�D�������U9��G��D��������4���Y����W	��C��\�ߊu�u�<�;�;�:����I����l ��Y�����0�
�4�
�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����T��Q1�����3�
�b�
�9�����&����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʲ�%�3�e�3�f�;�(��&����V ��R��E��������4���Y����W	��C��\�ߊu�u�<�;�;�:����I����l ��Y�����0� �;�e�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��h^��*ۊ� �f�l�4��8����H����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�
��(�D�������G��h\��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%��(߁�&¹��lU��h�����'�
�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����U9��Q1�����b�
�%�'�#�/�(���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����e�3�d�3��j�(�������]9��N��1��������}�D�������V�=N��U���;�9�2�%�1�m��������
9��h��Oʆ�����]�}�W�������lP��B�����d�d�&�'�0�o�E��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���3�'�0�d�g�.����K���5��h"��<������}�f�9� ���Y����F�D�����
�
� �3�%�8�G���
����lT��T��!�����
����_������\F��d��Uʦ�2�4�u�
��(�����֓�l��R	��@���u��
����2���+������Y��E��u�u�&�2�6�}�(ہ�����l��h_��*���
�c�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Q��R��*ۊ�
�
�0�
�`�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�����
�
�
�
��8�(��Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����7�3�0�
���(������� F��d:��9�������w�n�W������]ǻN�����9�%�m�7�1�8�(���&ù��A��_�Oʆ�������8���J�ƨ�D��^����u�<�;�9�'�e��������9��D1����l�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�A����U��R1��E���'�2�f�g�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������l^��B�����d�d�&�'�0�n�B��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������:�
�:�%�o�/���A����g"��x)��*�����}�u�8�3���B�����Y�����3�e�3�d�1��@ց�	����A��G1�����'�2�o����0���C���]ǻN�����9�4�
��1�0�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h��*���
�g�u�u���6��Y����Z��[N��*���
�1�
�b�w�}�8���8��ƹF��^	��ʴ�
�<�
�1��j�MϜ�6����l�N�����u�%�&�2�5�9�D��CӤ��#��d��Uʦ�2�4�u�%�$�:����M����q)��r/�����u�<�;�9�6���������\��x!��4��u�u�&�2�6�}��������lP��N��:����_�u�u�>�3�Ͽ�&����Q��_��U�����n�u�w�.����Y����Z��S
��E������]�}�WϽ�����]��r(�D��3�e�3�d��W�W������9F�N��U���6�>�o��w�	�(���0��ƹF�N�����!�o��u���8���B���F������!�o��u���8���B���F������u�u� �u���8���B���F������u�u� �u���8���B���F������,�o�����;���:���F�N��*���
�9�=�
�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y���Z��R�����u�u�����0���/����aF�N�����u�|�_�u�w�}�W���)����W9��N��U���
���
��	�%���Hӂ��]��G�U���u�u�<�
�2�����I����}F��s1��2������u�d�}�������9F�N��U���'�!�'�
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���Y�����E�����u�u� �u���8���&����|4�_�����:�e�n�u�w�}�WϿ�&����A��T�� ����
�����#���Q����\��XN�N���u�u�u�4��8����J����f2��c*��:���
�����l��������l�N��Uʴ�
�0� �;�c�g�8���*����|!��h8��!���}�d�1�"�#�}�^�ԜY���F��h�� ���`�o�����;���:����g)��]����!�u�|�_�w�}�W���	����	F��=��*����u�n�u�w�8�Ͻ�����]��=d�����_�u�u�'���(���&����_������;�u��l�f�e������ƹF��X�����}�u�u�u�w�<�(���Y����C9��\BךU���u�u�%�'�#�`�W�������F�N�����!�'�u�k�0�-�����ד�F9��1��*���'�y�u�u�w�}�������F��G1��E���d�3�
�b��-����U���F������u�k�2�%�1�m��������
9��h���ߊu�u�u�u�'�/����D�ƫ�C9��1��D���
�b�
�%�%�<��ԜY���F��h��*���=�
�u�k�0�-�����ד�F9��1��*���
�9�=�
�{�}�W���Yӏ��A��Z��F��u�'�
�
���(���J�ߓ�]9��Q1����_�u�u�u�w�3�'�������X��E��*ڊ�
�
� �f�n�4�(�������l�N��Uʼ�
�0�
�0�6�m�J�������9��1��*��
�;�'�3�5�)�(��Y���F��G1�����
�u�k�2�'�;�G���H���� Q��V�����;�e�_�u�w�}�W�������]9��
P�����
�
�
�
�"�n�N���&����A��d��U���u�4�
�0�"�3�E��Y����U9��Q1�����b�
�%�'�#�/�(��Y���F��G1�����
�u�k�2�'�;�G���H���� Q��V�����;�f�_�u�w�}�W�������]9��
P�����
�
�
�
�"�n�N���&����A��d��U���u�4�
�0�"�3�B��Y����U9��Q1�����b�
�%�'�#�/�(��Y���F��G1��U��2�%�3�e�1�l����Nʹ��l��dװ�ߊu�u�x�!�2�>����ӕ��G�V��&���8�u�3�!�2�.��������]�CךU���%��
�&��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F������u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�4������E�ƭ�l(��Q�����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӁ��l ��h��*���f�l�4�
�#�/�(���
����l�������%�:�0�&�w�p�W�������lV��h_�� ��l�4�
�!�%���������V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���'�
�
�
�����@����@��C1��*���'�
�0�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�g�3�8�f�}��������\��h��F���%�u�u�%�4�3����H���F��R ��U���u�u�u�u�w�}�W�������lV��h_�� ��l�4�
�!�%���������V�
N��*���&�
�:�<��f�W���Y���F�N�����u�}�%�6�9�)���������h��*���
� �f�l�6�����P�Ƹ�V�N��U���u�u�u�u�w�}�����֓�lW��B1�L���
�!�'�
�'�.�������F��h�����:�<�
�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����e�4�
�9��/�Ͽ�
����C��R��U���u�u�%�e�g�<�(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U´�
�<�
�1��e�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(߁�&����_��E��I���%�6�;�!�;�:���s���F�N��U���u�u�0�&�1�u��������lU�����ߊu�u�u�u�w�}�W���Y���F��1�����9�
�'�2�k�}�(߁�&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�m�G����ƭ�@�������{�x�_�u�w��(߁�����@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ڊ�
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F��	�֓�l��A��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(������O��_�����u�u�u�u�w�}�W���Y����9��R	��Hʥ�e�e�_�u�w�}�W���Y���V��^����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���F���*ۊ�%�#�1�%�2�}����Ӗ��P��N����u�
�
�
�'�+��������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��E���4�
�9�
�%�:�K���	����@��X	��*��u�u�u�u�w�}����s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��QN�����2�7�1�f�g�}����s���F�N��U���u�u�u�u�'�m�F���&����C��R�����:�&�
�:�>��L���Y���F�N��U���u�9�<�u�6���������F��R ��U���u�u�u�u�w�}�W���Y����lV��h�����%�0�u�h�'�m�F���&����9F�N��U���u�u�u�u�w�3�W���s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�
����������]F��X�����x�u�u�%�g�l����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��D���0�u�h�4��2�����ԓ�l�N��U���u�0�&�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]���%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�}��������]��[����h�4�
�!�%�t�^Ͽ��έ�l��D�����
�u�u�
���������G��d��U���u�u�u�u�w�}�WϮ�I�ד�A��S��*ڊ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1��*���
�'�2�4�$�:�W�������K��N�����4�
�9�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lW��G1�����0�u�h�4��2��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN�����:�&�
�:�>��W���	����F��R ךU���u�u�u�u�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y���F�N��U���
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W���Y���F��D��]���&�2�7�1�b�t����Y���F�N��U���u�u�u�u�w��(�������A��S��*ۊ�%�#�1�_�w�}�W���Y���F�N��ʼ�n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��1�����&�<�;�%�8�8����T�����h�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�%�f�-����DӇ��P	��C1��F؊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����R��[
��\ʡ�0�u�u�u�w�}�W���Y���F��h_�����i�u�
�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�g�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z �V�����1�
�m�|�#�8�W���Y���F�N��U���u�u�u�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���F�N�����3�}�%�&�0�?���PӒ��]FǻN��U���u�u�u�u�w�}�W���&����l��h����u�
�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����%�0�u�&�>�3�������KǻN��*؊�'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����	����[��G1�����9�f�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����}�%�6�;�#�1����I����C9��V��\���;�u�4�
�8�.�(�������F��1��*���|�|�!�0�w�}�W���Y���F�N��U���
�'�2�i�w��L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�`�e�6���������@��YN�����&�u�x�u�w�-�B�������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���<�u�4�
�>�����A����[��=N��U���u�u�u�u�w�}�W���Y����9��h��*���2�i�u�%�4�3��������l�N��U���u�u�u�u�w�8����Q����Z��S
��D���=�;�_�u�w�}�W���Y���F�N�����e�4�
�9��/���Y����9��h��N���u�u�u�u�w�}�W���YӃ����=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�L�֓�A��V�����'�6�&�{�z�W�W���&ƹ��C��h�����%�:�u�u�%�>����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�r�p�}����Y���F�N�����%�'�!�h�p�z�W������F�N��U���u�
�
�
�%�:�K���	����@��A]��E�ߊu�u�u�u�w�}����Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�;�!�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}�������F��SN�����;�!�9�2�4�l�JϮ�L�֓�C9��SG��U���;�_�u�u�w�}�W���Y���F��1�����u�h�%�`�g�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���
�
�
�%�!�9����Y����T��E�����x�_�u�u���(�������A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�`�d�4��1�(������R��X ��*���<�
�n�u�w�}�W���YӃ��Vl�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U���}�%�&�2�5�9�D��Y����l�N��U���u�u�u�u�w�}�WϮ�L�ד�C9��S1�����h�4�
�:�$�����&��ƹF�N��U���u�u�u�u�;�4�Wǿ�&����Q��^�����u�u�u�u�w�}�W���Y���F���*ۊ�%�#�1�%�2�}�JϮ�L�ד�C9��SUךU���u�u�u�u�w�}�W����ƥ�l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}�(ځ�&������^	�����0�&�u�x�w�}����H����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʥ�`�d�%�0�w�`��������_��h^�U���u�u�u�u�2�.�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�}�%�4�3��������[��G1�����0�
��&�f�;���Y������T�����2�6�e�h�6�����P����]�V�����
�:�<�
�w�}�(ځ�&����_�N�����u�u�u�u�w�}�W���Y����lS��h����u�
�
�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����<��'��8��(���&����R��P �����&�{�x�_�w�}�;���&����	��hV�����c�
�&�<�9�-����Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�^�����<�
�1�
�`�t����Y���F�N��U���u�u�u��;���������l��h]�U��<�
�<��%�����&¹��T9��UךU���u�u�u�u�w�}����Yۇ��@��U
��D��u�=�;�_�w�}�W���Y���F�N��*����'��:������O�����T�����g�e�_�u�w�}�W���Y���V��^�U���u�u�u�u�2�9���s���F�R ����u�u�0�1�'�2����s���K�V�����'�6�&�{�z�W�W�������@F��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���^�Ƹ�VǻN��U���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o����H�ƭ�WF��O�����
� �f�b�'�}�W�������l
��h^��\ʡ�0�_�u�u�w�}�W���Y�ƪ�l
��q��9���
�f�'�2�b�d�K���*����u	��{��*���3�
�e�
�d�W�W���Y���F�N��*����'��:��h����L���F��h��3����:�
�`�1��F߁�J���F�N��U���u�!�%�'�0�h�D��Y����U��W��D�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�E������F��R ךU���u�u�u�u�w�}�;���&����	��hV��*���
�`�u�h�>���������C9��1��*��
�g�_�u�w�}�W���Y����Z ��N��U���0�1�<�n�w�}����	����@��=N��U���4�&�2�u�%�>���T���F��X�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������A��N���ߊu�u�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�Փ�@��N��ʻ�!�}�%�6�9�)���������h��*���
� �f�l�6�����P����[��N��U���u�u�u�u�'�i��������9��D1����f�i�u�
��(����H����lT��B1�M���n�u�u�u�w�}�W���YӖ��l��Q�����d�&�'�2�e�m�K���&ǹ��U ��h_��*ڊ�
� �a�d�'�f�W���Y���F�N��*ފ� �3�'�0�f�m��������Z�G1�����0�
�
�
�����K����9F�N��U���u�u�u�
��(�����ד�l��R	��C���h�%�a�7�1�8�(ށ�&¹��U��[��F�ߊu�u�u�u�w�}�W���&Ź��U ��h��*ڊ�
�0�
�`�w�`��������A9��R1��G���
�b�
�f�]�}�W���Y���F�G1�����0�
�
�
������J�����h�����d�0�e�d�1��Aց�J���F�N��U���u�%�c�7�1�8�(���&ù��A��\�I���
�
� �3�%�l����K����_��G]�U���u�u�u�u�w�}��������A9��1�����2�g�g�i�w��(�������l��h_�� ��f�%�n�u�w�}�W���Y�����h�����0�e�e�&�%�:�D��E�Ƽ�9��Q��*ۊ�
�
�
� �c�j���Y���F�N��U���
�
� �3�%�8�G���
����lU��R�����7�3�0�
���(݁�����l��=N��U���u�u�u�u�w��(�������lW��h�����a�u�h�%�o�?����&¹��9��Q��Dۊ�f�_�u�u�w�}�W���Y�Ƽ�9��Q��*���
�
�
�0��h�W��	�ޓ�F ��E1�����g�3�
�d��n�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�#�8����Y����VF��G1��*���|�:�u�=�w�)��������VH�d��Uʴ�
��3�8�6�.���������T��U´�
��3�8�w�-�������T9��S1�A���-�!�:�1��(�D���	����A��h^��*ۊ� �f�l�4��2��ԜY�Ʈ�T��N��U���6�&�u�%������
���F�N��U���;�4�
��$�l����I���9F�N��U���u�u�u�3��u��������\��h_��U���6�|�4�1�9�)��������W9��G��U���;�u�u�u�w�}�W���Y�����y=�����h�4�
��$�o����H���F�N��U���u�0�&�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�u�u�9�}��ԜY���F�N�����%��
�!��.�(���G���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�:��8�����Փ�F9�� 1��U���%�6�;�!�;�l�G���PӒ��]l�N��U���u�u�u�u�w�<�(������F��h=�����3�8�e�_�w�}�W���Y���F��DךU���u�u�u�u�w�}�W���	����U��S�����
�!�
�&��f�W���Y���F�N�����3�_�u�u�w�}�W�������C9��h��*���
�u�k�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]´�
�:�&�
�8�4�(���Y����U9��Q1�����b�
�%�1�9�t�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W���Y����_��N��U���u�u�u�u�w�}����*����Z�V��!���f�3�8�g�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����A�	N��U���u�u�u�u�w�}����*����Z�6��W�ߊu�u�u�u�9�}����s���V��G�����_�u�u�x�w�-����Y����T��E�����x�_�u�u�'�9����
����l��TN����0�&�4�
�2�}��������B9��h��*���
�y�0�<�4�3�D���&����CT�N�����;�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$�������^9����U���}�0�<�6�9�n����AĹ��[��G1�����9�d�e�|�~�)����Y���F�N�����;�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����\��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h��ʴ�&�2�u�'�4�.�Y��s���R��S�����2�
�'�6�m�-����
ۇ��@��CB�����2�6�0�
��.�F������F�U�����u�u�u�<�w�u��������]��[����h�4�
�!�%�t�W���Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\���=�;�_�u�w�}�W���Y����W
��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��9���Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������R��P �����&�{�x�_�w�}��������@��Y1�����u�'�6�&��-�������T9��R��!���g�3�8�d�w�%��������lU��h����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GT��D��\ʴ�1�;�!�}�/�)����&����Q��N�����:�&�
�#��t�^������F�N��U���4�
�0�1�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���&�2�7�1�f�i�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4��)���	�֓�l��A�����<�y�%�e�f�<�(���&����Z�G1�����9�
�;�&�0�}�(݁�	����l��D��U���
�
�%�#�3�4�(���UӖ��lW��G1�����
�<�|�u�w�?����Y���F�N��U���%�&�2�7�3�l�C��Y�μ�9��h��*���&�2�h�4��2��������O��EN��*ۊ�%�#�1�<��4�W���	����@��X	��*���:�u�%�`�g�<�(���&����Z������!�9�2�6�g�}����&ƹ��R��[
�����2�h�4�
�8�.�(�������	����*ڊ�%�#�1�<��4�W���	����@��X	��*���:�u�%�e�f�<�(���&����Z������!�9�2�6�g�}����	����A������!�9�2�6�g�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����l��F1��*���
�&�
�y�6���������OǻN�����_�u�u�u�w�}�W���Y����Z��S
��G���h�}�4�
�8�.�(�������F��h��*���$��
�!��.�(�������\��G1�����1�d�a�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h_�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�d�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h_�U��}�%�6�;�#�1�F��DӇ��p5��D��U���;�:�g�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u��������B9��h��*���
�y�2�%�1�m��������
9��h
���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�b�u�j�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����4�
�:�&��2����Y�ƫ�C9��1��D���
�b�
�%�3�3�^���s���V��G�����_�_�u�u�z�<�(���&����_��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��W�����;�%�:�u�w�/����Q����`9��ZGךU���0�<�_�u�w�}�W���Y���R��^	�����l�i�u�4������Iӂ��]��G��U���6�;�!�9�f�l�L���YӃ����T��N�ߠu�u�x�u�'�.��������R��P �����&�{�x�_�w�}��������lU��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�f�u�h��<�(���
����T��N�����e�4�
�9�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�n�u�u�2�9��������9l�N�U���&�2�7�1�d�m�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4��4�(�������@��Q��D���-�!�:�1��(�D���	��ƹF��R	�����u�u�u�u�w�}�W���
����W��^��H���4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�������V��T��F���
�m�
�g�j�<�(���
����9��G�U���0�1�%�:�2�.�}�ԜY�����D�����a�u�&�<�9�-����
���9F������7�1�a�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
�
�%�!�9�}���Y����]l�N��U���u�u�u�4��4�(���&���F��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
��-����P���F��SN�����&�_�_�u�w�p��������W9�������%�:�0�&�w�p�W�������T9��S1�*���<�;�%�:�w�}����
�έ�l��E����<�
�&�$���ށ�
������h�����_�u�u�0�>�W�W���Y���F�N��*���
�1�
�`�k�}����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�4�
�:�$�����&���R��C��\���4�1�}�%�4�3��������[��h_�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��i�����Ƽ�\��D@��X���u�4�
�<��9�(�������]9��X��U���6�&�}�%�$�<����	����l��F1��*���
�&�
�y�'�o������ƹF��R	�����u�u�u�u�w�}�W���
����W��N�U»�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�E���&����]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��Dʴ�&�2�u�'�4�.�Y��s���R��^	�����d�4�&�2��/���	����@��G1�����u�%�&�2�4�8�(���
�ד�@��N��@���4�
�9�|�w�}�������F�N��U���u�%�&�2�5�9�O���D�΢�GN�V�����
�:�<�
�w�}��������B9��h��*���
�|�4�1��-��������Z��S�����4�!�|�u�9�}��������_	��T1�Hʥ�`�e�4�
�;�t�L���YӃ����T��N�ߠu�u�x�u�'�.��������R��P �����&�{�x�_�w�}��������l_��V�����'�6�o�%�8�8�ǿ�&����GJ��G1�����0�
��&�f�;���Y����9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�l�u�h��2�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N�����%�6�;�!�;�:���DӇ��@��CG��U���u�4�
�:�$�����&���C9��1��*���|�n�u�u�2�9��������9l�N�U���&�2�6�0��	����������^	�����0�&�u�x�w�}��������V��c1��D���8�e�4�&�0�����CӖ��P�������7�1�d�|�w�}�������F���]���&�2�7�1�f�t����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����l ��h^��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�o����HӇ��Z��G�����u�x�u�u�6�����
����g9��1�����4�&�2�
�%�>�MϮ�������D�����d�c�_�u�w�8��ԜY���F��F��*���
�1�
�a�~�)����Y���F�N�����2�6�0�
��.�E������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�&�2�4�8�(���
�ԓ�@��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����0�
��&�d�;�������]F��X�����x�u�u�4��4�(�������@��Q��G���&�2�
�'�4�g��������C9��P1����c�_�u�u�2�4�}���Y���Z �V�����1�
�c�|�#�8�W���Y���F������6�0�
��$�n����K���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�&�2�6�2��#���J����lT�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}���YӃ��G��S]�� ��b�%�u�h�u�� ���Yۏ��_��X�����m�'�2�f�o�`��������_��G�����w�w�_�u�w���������\��1��*��
�f�i�u�w�}�W���	�֓�l��D�����u�!�%�3��d�(��I���W����ߊu�u�u�u���(���
����F�Q=�����'��:�
�b�;�(��&���FǻN��U���
�
�
�;�$�:� ���Yے��l ��W�����|�h�r�r�w�1��ԜY���F��1�����<�n�_�u�w�p�����֓�lW��B1�L���
�0�4�&�0�}����
���l�N�����e�3�d�3��j�(�������@��h����%�:�0�&�6�����	����l��F1��*���
�&�
�y�6�����
����g9��1����_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��G1�����9�2�6�d�j�<�(���&����l5��D�����d�u�'�}�'�>��������lW������6�0�
��$�n����K�����YNךU���u�u�u�u�%��(߁�&¹��lU��h�����h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���&����U9��Q��Bӊ�%�6�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���'�
�
�
�����@����@��CN�U���
�
�
�
��(�D�������R��V�����
�0�n�u�w�:����I����l ��Y�����0�<�1�a�k�}�(݁�����l�N�����e�3�d�3��j�(�������_��h_��Hʳ�
�!��'��2�(�������_��N�����3�e�3�d�1��@ց�����l��V1�I����9�
�:��2���&����^��=N��U���
�
�
�
��(�D�������U9��O1�I���
�
�;�&�0�W�W���5����u	��{��*Ҋ�
� �f�f�'�}�Jϭ�����Z��R�� �&�2�0�}��1�(���&����l^��R	��C���~� �&�2�2�u��������ET��G����u�x�%�e�g�<�(���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�I�֓�C9��S1��*���
�&�<�;�'�2�W�������@N��1�����9�y�%�e�g�<�(���&����l�N�����u�u�u�u�>�}�_�������l
��^��U���
�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�
�%�!�9���������h^�����1�_�u�u�w�}����s���F�N�����e�4�
�9��3����E�Ƽ�9��V�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���&ù��Z��^	�����;�%�:�0�$�}�Z���YӖ��lV��Y1�����&�2�
�'�4�g��������lV��N��E���%�0�y�%�g�m������ƹF��R	�����u�u�u�3��<�(���
����T��N�����e�4�
�9�~�}����s���F�N�����e�<�
�<�w�`����I���F�N�����u�u�u�u�w�}����I����@��S��*ڊ�
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����9��h��*���&�2�4�&�0�}����
���l�N��E���4�
�9�
�9�.����
����C��T�����&�}�
�
��-����Y����9��h��*���2�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����H����E
��N�����u�u�u�u�w�}����H����E
��^ �����h�%�e�d�6����Y���F��[�����u�u�u�u�w��(ށ�	����l��D��I���
�
�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ڊ�
�;�&�2�6�.��������@H�d��Uʥ�e�d�<�
�>���������PF��G�����%�e�d�u���(����Ƽ�9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(ށ�	����O��_�����u�u�u�u�w��(ށ�����Z�G1��D�ߊu�u�u�u�;�8�}���Y���F�G1��D���
�<�u�h�'�m�F�����ƹF�N�����3�u�u�u�2�9��������9l�N�U���
�%�#�1�>�����
������T��[���_�u�u�
��-��������T9��D��*���6�o�%�:�2�.��������WJ��h_�����1�%�0�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����R��[
��U���;�_�u�u�w�}�W���&¹��l��h�����i�u�
�
�'�+��ԜY���F��D��U���u�u�u�u�'�l��������l��R�����4�
�9�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��1��*���u�&�<�;�'�2����Y��ƹF��h_�����2�4�&�2��/���	����@��h_����%�0�y�%�f�<�(���P�����^ ךU���u�u�3�}�6�����&����P9��
N��D���
�9�|�u�?�3�}���Y���F�G1�����<�u�h�%�f�W�W���Y�Ʃ�@�N��U���u�u�%�d�>�����DӖ��l��PUךU���u�u�;�u�1�}�W�������A	��D����u�x�u�
��-��������TF��D��U���6�&�{�x�]�}�W���&����_��Y1�����&�2�
�'�4�g��������lT��G1�����
�
�%�#�3�-����Y����V��=N��U���u�3�}�4��2��������F�G1�����9�|�u�=�9�W�W���Y���F��1��*���
�;�&�2�k�}�(݁�	����l�N��Uʰ�&�u�u�u�w�}�W���	�ԓ�C9��S1��*���u�h�%�g�6���������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�g�<�
�<�w�.����	����@�CךU���
�
�;�&�0�<����&����\��E�����
�y�%�g�'�8�[Ϯ�K����E
��=N��U���<�_�u�u�w�}��������]��[����h�%�g�4��1�^������F�N��U���%�g�<�
�>�}�JϮ�K���F�N�����u�u�u�u�w�}��������TF���*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w��(߁�&�����h�����0�e�e�&�%�:�D��s���K�G1��E���e�4�
�9�w�.����	����@�CךU���
�
�
�
��-��������]9��X��U���6�&�}�%�4�q��������V��c1��G���8�d�u�-�#�2�܁�����l��=N��U���<�_�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�ԓ�@��N��ʻ�!�}�-�!�8�9�(���J�ѓ�F�V�����
�#�
�|�~�}����s���F�N�����e�0�e�4��1�W������]��[����_�u�u�u�w�1��ԜY���F�N��A���0�e�4�
�;�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�
���(���DӖ��l��Q�����e�&�'�2�e�j�}���Y���C9��1��D���
�9�u�&�>�3�������KǻN��*ފ�
�
�
�%�!�9��������\������}�%�6�y�6�����
����g9��1����u�-�!�:�3����N����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������F��SN�����-�!�:�1��(�D���	���R��X ��*���
�|�|�u�?�3�}���Y���F�G1��E���d�4�
�9�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��1�����4�
�9�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�
�
�
��}�JϮ�M����U��R1��D���'�2�g�e�]�}�W��Y����9��1��*���u�&�<�;�'�2����Y��ƹF��hZ��*���
�%�#�1�6�.���������T��]���6�y�4�
�>�����*����9��Z1�U���!�:�1�
�"�n�@���P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o����H�ƭ�WF��CF�����:�1�
� �d�j����Y����\��h��*���|�u�=�;�]�}�W���Y���C9��1��E���
�9�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��R1�����9�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=N��U���
�
�
�u�j�-�C�������V9��1�����g�a�_�u�w�p�W���&¹��9��h��U���<�;�%�:�2�.�W��Y����lR��h��*���#�1�4�&�0�����CӖ��P�������4�
�<�
�$�,�$�������^9�������1�
� �f�`�-�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�g�1�0�F����Ƣ�GN��O�����
� �f�b�'�}�W�������l
��h^��\���=�;�_�u�w�}�W���Y����9��1��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���&ǹ��V9��V�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9F���*���3�'�d�0�g�l����M¹��Z�=N��U���u�'�
�
���(���J�ߓ�C9��C��*���=�;�}�8��8�(��Q���A��N�����u�u�u�u�'�i��������9��D1����e�_�u�u�������ד�lV��h��A���%�u�h�_�w�}�W���&ǹ��U ��h��*ڊ�
�0�
�e�w�5��������T9��F�U���d�|�0�&�w�}�W���YӁ��l ��h��*���f�l�4�
�2�(���s���C9��U�����
�
�
�
�"�i�B���Y���F�N�����3�e�3�d�1��@ց�	����F��N�����!�%�'�2�b�n�G���Y�����RNךU���u�u�
�
�"�;����H�ד�l��h\�N���u�%�a�7�1�8�(ށ�&¹��U��\��F��u�u�u�u�w�-�C�������V9��1�����g�b�"�0�w�)��������V�
N��R���9�0�_�u�w�}�W���&����U9��Q��Bӊ�%�'�!�'��f�}���Y����lS��h�����<�
�<�u�$�4�Ϯ�����F�=N��U���
�
�%�#�3�4�(���&����T��E��Oʥ�:�0�&�%�b�m��������lS��h�����%�0�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&ƹ��R��[
��U���;�_�u�u�w�}�W���&ƹ��R��[
�����2�i�u�
���������F�N�����u�u�u�u�w�}����I����E
��^ �����h�%�`�e�6���������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʥ�`�e�<�
�>�}����Ӗ��P��N����u�
�
�
�9�.����
����C��T�����&�}�
�
�{�-�B���	������h^�����1�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����I����E
��N�����u�u�u�u�w�}����I����@��S��*ߊ�n�u�u�u�w�8����Y���F�N��*ߊ�
�;�&�2�k�}�(ځ�&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�`�d�4��1�(���
����@��YN�����&�u�x�u�w�-�B�������W9��h��*���<�;�%�:�w�}����
�μ�9��V�����%�`�d�4��1�(������F��P��U���u�u�<�u��-��������Z��S��*ߊ�
�%�#�1�~�)����Y���F�N��*ߊ�
�%�#�1�>�����DӖ��lW��G1���ߊu�u�u�u�;�8�}���Y���F�G1��D���
�9�
�;�$�:�K���&ƹ��R��[
�����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}�(ځ�&����Z��D��ʥ�:�0�&�u�z�}�WϮ�L�ד�]9��P1�����
�'�6�o�'�2����	�ӓ�F��1�����y�%�`�d�6�����Y����V��=N��U���u�3�}�4��2��������F�G1��D���
�9�|�u�?�3�}���Y���F�G1��D���
�<�u�h�'�h�F�ԜY���F��D��U���u�u�u�u�'�h�F���&����[��h[��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w��(߁�&�����h�����0�e�e�&�%�:�E��s���K�G1��E���e�4�
�9�w�.����	����@�CךU���
�
�
�
��-��������]9��X��U���6�&�}�%�4�q��������V��c1��G���8�d�u�-�#�2�܁�����l��=N��U���<�_�u�u�w�}����Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
�ԓ�@��N��ʻ�!�}�-�!�8�9�(���J�ѓ�F�V�����
�#�
�|�~�}����s���F�N�����e�0�e�4��1�W������]��[����_�u�u�u�w�1��ԜY���F�N��C���0�e�4�
�;�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�
���(���DӖ��l��Q�����e�&�'�2�e�h�}���Y���C9��1��D���
�9�u�&�>�3�������KǻN��*܊�
�
�
�%�!�9��������\������}�%�6�y�6�����
����g9��1����u�-�!�:�3����N����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������F��SN�����-�!�:�1��(�D���	���R��X ��*���
�|�|�u�?�3�}���Y���F�G1��E���d�4�
�9�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��1�����4�
�9�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�
�
�
��}�JϮ�O����U��R1��D���'�2�g�m�]�}�W��Y����9��1��*���u�&�<�;�'�2����Y��ƹF��hX��*���
�%�#�1�6�.���������T��]���6�y�4�
�>�����*����9��Z1�U���!�:�1�
�"�n�@���P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o����H�ƭ�WF��CF�����:�1�
� �d�j����Y����\��h��*���|�u�=�;�]�}�W���Y���C9��1��E���
�9�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��R1�����9�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=N��U���
�
�
�u�j�-�A�������V9��1�����g�g�_�u�w�p�W���&¹��9��h��U���<�;�%�:�2�.�W��Y����lP��h��*���#�1�4�&�0�����CӖ��P�������4�
�<�
�$�,�$�������^9�������1�
� �f�`�-�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�g�1�0�F����Ƣ�GN��O�����
� �f�b�'�}�W�������l
��h^��\���=�;�_�u�w�}�W���Y����9��1��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���&Ź��V9��V�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9F���*���3�'�d�0�g�l����Oʹ��Z�=N��U���u�'�
�
���(���J�ߓ�C9��C��*���=�;�}�8��8�(��Q���A��N�����u�u�u�u�'�k��������9��D1����m�_�u�u�������ד�lV��h��A���%�u�h�_�w�}�W���&Ź��U ��h��*ڊ�
�0�
�`�w�5��������T9��F�U���d�|�0�&�w�}�W���YӁ��l ��h��*���f�l�4�
�2�(���s���C9��U�����
�
�
�
�"�i�D���Y���F�N�����3�e�3�d�1��@ց�	����F��N�����!�%�'�2�b�n�G���Y�����RNךU���u�u�
�
�"�;����H�ד�l��h\�N���u�%�c�7�1�8�(ށ�&¹��U��^��F��u�u�u�u�w�-�A�������V9��1�����g�`�"�0�w�)��������V�
N��R���9�0�_�u�w�}�W���&����U9��Q��Bӊ�%�'�!�'��f�W���	�ޓ�l��R�����7�3�0�
���(�������]ǑN��X���
�
�
�
��-��������]F��X�����x�u�u�%�o�m��������W9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�
�&��q��������l ��V�����u�u�7�2�9�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1����u�;�u�:��8�����Փ�F9�� 1��U���%�6�;�!�;�l�G���PӒ��]FǻN��U���u�u�
�
���(������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�
�
�
���������R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}����I����Z�G1�����0�
�
�
������M��ƓF�C��*Ҋ�
�
�
�%�!�9�����Ƽ�\��D@��X���u�%�m�e�2�l��������@��h����%�:�0�&�6�����	����l��F1��*���
�&�
�y�2�4����J���� ^��G\��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�:�}�0�>�>��������9��S�����;�!�9�d�g�t�^Ϫ���ƹF�N��U���
�
�
�
��-����E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���
�
�
�
�'�+���Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�'�e�F���I���C9��U�����
�
�
�
�2��E��s���K��hV��*���
�%�#�1�6�.��������@H�d��Uʥ�m�d�0�e�6�����
����l��TN����0�&�4�
�2�}��������B9��h��*���
�y�0�<�4�3�D���&����CT�N�����;�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$�������^9����U���}�0�<�6�9�n����AĹ��[��G1�����9�d�e�|�~�)����Y���F�N��*Ҋ�
�
�
�%�!�9�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F���*ۊ�
�
�%�#�3�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠu�u�%�m�f�8�F��Y����Q��R��*ۊ�
�
�0�
�b�f�}���Y����l^��h��*���#�1�4�&�0�}����
���l�N��M���0�d�4�
�;���������PF��G�����4�
�0�u�'�.��������l��h��*���0�<�6�;�d�;�(��&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$���݁�
������ ��]°�<�6�;�f�1��O؁�K����C9��Y�����e�|�|�!�2�}�W���Y���F��hV��*���
�%�#�1�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����h_��*ۊ�%�#�1�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���%�m�7�3�2��(���&¹��lR��h�I���u�u�u�u�'�e��������9��D1����c�"�0�u�#�-����L���F�_��U���0�_�u�u�w�}����&ù��9��h]�*���'�!�'�
�l�}�WϮ�A����U��1��E���3�
�e�
�d�a�W���Y�����h��*���
� �f�l�6���������[����*���
�c�}�|�j�z�P������F�N�����7�3�0�
���(�������
]ǻN��*Ҋ� �3�'�d�2�l�F���&����CU�
NךU���u�u�
�
�"�;����H�֓�l��h]�U���;�}�8�
�2��A���P���A�R��U���u�u�u�2�'�;�G���H���� Q��V�����;�`�_�u�w��(�������l��h\�� ���m�%�u�h�]�}�W���Y����U9��Q1�����b�
�%�'�#�/�(������G��E��@��e�u�u�d�~�8����Y���F��hV�� ���'�0�d�d�$�/���L���F��G1��*��
�d�i�u��1�(���&����l^��R	��C���u�u�u�:�9�2�G������V��d