-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��LӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�c��b�b��}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e�o��u���8���&����|4�_�����:�e�n�u�w�<�(���Cӯ��`2��{!��6�ߊu�u�
�
�'�+���0�Ɵ�w9��p'�����u�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���&����_�'��&������_�w�}�(���Y����g"��x)��*�����}�d�3�*����P���F��1��*���u�u�����0���s���C9��R1�Oʚ�������!���6���F��@ ��U���_�u�u�
���(������)��=��*����n�u�u�'�i���Cө��5��h"��<������}�f�9� ���Y����F�G1�����4�
�9�u�w��W���&����p]ǻN��*���u������4���:����U��S�����|�_�u�u����������}F��s1��2���_�u�u�
���W���,�Ɵ�w9��p'��#����u�f�u�8�3���B�����h��*���#�1�o����3���>����F�G1����o������0���/����aF�N�����u�|�_�u�w��(���&����_�!��U���
���n�w�}�������)��=��*����
����u�FϺ�����O��N�����0�e�4�
�;�}�W���Y����)��tUךU���
�
�
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ޓ�lW��G1����������4�ԜY�Ƽ�S�!��U���
���
��	�%���Y����G	�UךU���
�`�4�
�;�}�W���Y����)��tN����n�_�4�6�>�8����Y����EF����1��m�3�e�<�w�}�WϿ�����G��x<��2������
���Mύ�+����9F������!�u�����%���6����u)��QN�����o�4�6�<�2�)����
���D��*��B���
�y�9�
�'�o�Fځ�U����l/��b:��,���6�-�����#���6���.��h'�� �����h�y���9���&������M^����m�x�y����"���5����S�^�EƝ�������J�������5��n ��9���h�d�m�m�g�q�;��� ����g[��&��*���
��h�:�2��$���7����S��{=��,����h�y����(���H����{*��d7��9���b�`�(�n�w�}��������R��X ��*���<�
�u�u���8���Y���A��N�����!�;�u�%�4�3��������\��c*��:���u�h�r�r�]�}�W���
������d:��ۊ�&�
�u�u���8���&����|4�W�����:�e�u�h�u�m�G��I����V��^�W�ߊu�u�:�&�6�)����-����l ��h_��U���
���
��	�%���@ӂ��]��G��H���e�e�e�e�g�m�G��I���9F������!�4�
��$�n����K����g"��x)��*�����}�l�3�*����P���V��^�E��e�e�e�d�g�f�W�������R��V��!���a�3�8�f�m��3���>����v%��eN��Lʱ�"�!�u�|�m�}�G��I����V��^�E��n�u�u�6�9�)����	����@��Q��A��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����D��N�����!�;�u�%���ف�
����	F��s1��2������u�f�}�������	[�^�E��e�e�e�d�g�m�U�ԜY�Ư�]��Y�����
�!�
�&��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�w�_�u�w�2����Ӈ��`2��CV�����u�u��
���(���-���_��X����u�h�w�e�g�m�G��I����V��UךU���:�&�4�!�6��#���@����l^�=��*����
����u�NϺ�����O�
N��E��e�e�e�d�g�m�G��B�����D��ʴ�
��&�d��.�(���Y����)��t1��6���u�d�u�:�9�2�G���D����V��^�D��e�e�e�w�]�}�W���
������d:�����3�8�d�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E���_�u�u�:�$�<�Ͽ�&����GW��Q��D���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V�=N��U���&�4�!�4��	���&����T�=��*����
����u�NϺ�����O�
N��E��e�d�e�e�g�m�G��B�����D��ʴ�
��&�d��.�(��Cӵ��l*��~-��0����}�l�1� �)�W���C���V��_�E��e�e�e�e�l�}�WϽ�����GF��h=����
�&�
�a�m��3���>����v%��eN��Lʱ�"�!�u�|�m�}�G��I����V��^�E��n�u�u�6�9�)����	����@��h��*���o������!���6���
F��@ ��U���o�u�e�e�f�m�G��I����V��d��Uʶ�;�!�;�u�'��(���N����lW��N��1��������}�F�������V�S��E��e�e�e�e�g�m�G��[���F��Y�����%��
�!�o�;���Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�e�e�u�W�W�������]��G1��*���l�3�8�d�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�E��w�_�u�u�8�.��������l��1����u�u��
���(���-���_��X����u�h�w�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lV�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
����9��N��1��������}�GϺ�����O�
N��W�ߊu�u�:�&�6�)��������_��hX��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�D���_�u�u�:�$�<�Ͽ�&����G9��\��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[�*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��d�e�w�_�w�}��������C9��Y����
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�d�d�w�]�}�W���
������T�����f�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�d�d�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�d�g��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�f�m�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�l�F���s���P	��C��U���6�;�!�9�d��G��*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�F��I��ƹF��X �����4�
�:�&��+�(���Y����)��t1��6���u�e�1�"�#�}�^��Y���9F������!�4�
�:�$�����H����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����K���5��h"��<������}�w�2����I����D��UךU���:�&�4�!�6�����&����lW��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}��������EP��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��h_��U���
���
��	�%���Jӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�D��u�u�6�;�#�3�W�������l
��1��Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�D��n�u�u�6�9�)����	����@��AX��G��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[�*��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�d�n�u�w�>�����ƭ�l��D�����d�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�d�d�w�]�}�W���
������T�����f�
��o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�d�d�f�f�W�������R��V�����
�#�g�f�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�d�g�m�U�ԜY�Ư�]��Y�����;�!�9�f���Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�l�F��B�����D��ʴ�
�:�&�
�!�o�4��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��n�u�u�6�9�)����	����@��AX��E��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��n�u�u�6�9�)����	����@��A_��A��o������!���6���F��@ ��U���o�u�e�e�g�l�G��[���F��Y�����%�6�;�!�;�l�(��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�D��n�u�u�6�9�)����	����@��A_��G��������4���Y����W	��C��\��u�e�e�e�g�m�F���s���P	��C��U���6�;�!�9�f��W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�W�ߊu�u�:�&�6�)��������_��h_��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�:�$�<�Ͽ�&����G9��_��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�`��}�W���&����p9��t:��U���u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D�����d�u�u����>���<����N��
�����e�u�h�w�g�m�G��I���9F������!�4�
�:�$�����?���5��h"��<������}�f�9� ���Y���F�_�D��e�e�n�u�w�>�����ƭ�l��D�����f�u�u����>���<����N��
�����e�u�h�w�g�m�G��H���9F������!�4�
�:�$�����H����`2��{!��6�����u�d�w�2����I����D��^�E��d�w�_�u�w�2����Ӈ��P	��C1��DҊ���u�u���8���&����|4�Y�����:�e�u�h�u�l�F��H����W��_�����u�:�&�4�#�<�(���
����^��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��B�����D��ʴ�
�:�&�
�!�o�1���Cӵ��l*��~-��0����}�d�1� �)�W���C���W��_�D��n�u�u�6�9�)����	����@��A_��D���u��
����2���+������Y��E���h�w�e�e�g�l�G��B�����D��ʴ�
�:�&�
�!�o�1���Cӵ��l*��~-��0����}�d�1� �)�W���C���W��_�D��n�u�u�6�9�)����	����@��A_��F���u��
����2���+������Y��E���h�w�e�e�g�l�F��B�����D��ʴ�
�:�&�
�!��B��*����|!��h8��!���}�u�:�;�8�m�W��[����W�=N��U���&�4�!�4��2����Ź��	F��s1��2������u�b�9� ���Y���F�^�E��u�u�6�;�#�3�W�������l
��1��3�������w�}�#���6����e#��x<��@���:�;�:�e�w�`�U��H����W��_�D��d�d�d�d�f�l�F��H����W��_�D��d�n�u�u�4�3����Y����\��h��G��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��d�e�n�u�w�>�����ƭ�l��D��Ҋ�u�u��
���(���-���F��@ ��U���o�u�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�d��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��_�����u�:�&�4�#�<�(���
����T��r/��U���
���
��	�%���Hӂ��]��G��H���d�d�d�e�g�m�L���YӅ��@��CN��*���&�
�#�g�f�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����W��^�����u�:�&�4�#�<�(���
����R��q(��3��������4���Y����W	��C��\��u�d�d�d�f�l�F��H����W��L�U���6�;�!�;�w�-��������9��N��1��������}�E�������V�S��E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)���&����	F��s1��2������u�f�}�������	[�_�D��d�e�w�_�w�}��������C9��Y����
�b�o����0���/����aF�N�����u�|�o�u�g�m�G��I����l�N�����;�u�%�6�9�)���&����	F��s1��2������u�f�}�������	[�_�D��d�e�w�_�w�}��������C9��Y����
�b�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�d�d�d�l�}�WϽ�����GF��h�����#�m�d���g�$���5����l0��c!��]��1�"�!�u�~�g�W��H����W��_�D��n�u�u�6�9�)����	����@��A_��G��e�o�����4���:����W��S�����|�o�u�d�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>�������� ��q(��U���
���
��	�%���Jӂ��]��G��H���d�d�d�d�f�l�F��H����W�=N��U���&�4�!�4��2�����ғ�V��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lT��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����W��^�N���u�6�;�!�9�}��������E_��T��!�����
����_�������V�S��E��e�e�e�n�w�}��������R��X ��*���
�u�u����>���<����N��S�����|�o�u�d�f�f�W�������R��V�����
�#�
�u�w�	�(���0����p2��F����!�u�|�o�w�l�G��Y����\��V �����:�&�
�#��}�W���&����p9��t:��U��1�"�!�u�~�g�W��H��ƹF��X �����4�
�:�&��+�B��Cӵ��l*��~-��0����}�a�1� �)�W���C���V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�f�f�g�$���5����l0��c!��]���:�;�:�e�w�`�U��[���F��Y�����%�6�;�!�;�n�C��*����|!��h8��!���}�u�:�;�8�m�W��[����l�N�����;�u�%�6�9�)����K����g"��x)��*�����}�u�8�3���Y���W��d��Uʶ�;�!�;�u�'�>�����Փ�\��c*��:���
�����}�������	[�_�N���u�6�;�!�9�}��������EU��V��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��_�E���_�u�u�:�$�<�Ͽ�&����G9��\��C��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�D��e�n�u�u�4�3����Y����\��h��G��u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��Y����
�`�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�d�d�d�l�}�WϽ�����GF��h�����#�g�f�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�d�e�f��}���Y����G�������!�9�f�
�`�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�f�l�F��Y����\��V �����:�&�
�#��}�W���&����p9��t:��U��1�"�!�u�~�g�W��[���F��Y�����%�6�;�!�;�n�G��*����|!��h8��!���}�u�:�;�8�m�W��[����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�g�w�2����I����D��^�E��e�e�e�e�g�m�L���YӅ��@��CN��*���&�
�#�g�`��1���Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���W��_�D��d�d�d�d�f�l�F��H����l�N�����;�u�%�6�9�)���&����V��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��N�&���������W������\F��T��W��n�u�u�6�9�)����	����@��A]��E��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[�*����o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��d�e�d�d�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�f��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�l�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s�����Y������3�8�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��^�D��u�u�4�!�>�(�ϸ�����\��PN����;�n�u�u�6�)����Ӏ��l��X
��ʺ�u�%��
�$�}�W�������@F��X ��N���u�&�2�4�w�-��������`2��C_�����u�u��
���L���Yӕ��]��V�����1�
�c�o���2���s���@��V��*ڊ�;�&�2�o���;���:����g)��]����!�u�|�_�w�}����Ӗ��l��PN�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��u�u�&�2�6�}�(߁�	����l��D��Oʆ�����]�}�W�������lV��G1�����0�u�u����>���D����l�N�����u�
�
�;�$�:�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��h_�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�.����Y����R��[
�����2�o�����4�ԜY�ƿ�T����*���#�1�%�0�w�}�#���6����	[�I�U���&�2�4�u����������g"��x)��*�����}�d�3�*����P���F��P ��U���
�'�2�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�f�W���
����_F��1��*���
�;�&�2�m��3���>����F�D�����
�
�%�#�3�-����Y����)��tN�U��n�u�u�&�0�<�W���&����Z�=��*����
����u�FϺ�����O��N�����4�u�
�
�%�:�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��B�����Y�����4�
�9�
�9�.���*����|!��d��Uʦ�2�4�u�
��-����	����	F��s1��2���o�u�e�n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��G1�L���2�f�l�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӂ��l ��Y�����u��
����2���+������Y��E��u�u�&�2�6�}�$���0����G9��1����l�u�u����>���<����N��
�����e�n�u�u�$�:����	����l��F1��*���
�&�
�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�1��o�W���6����}]ǻN�����9�2�%�3��j�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��&����,� �
�f�����A���5��h"��<������}�f�9� ���Y����F�D�����&�0�
�0��e�O��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��V�����&�$��
�#�����Y�Ɵ�w9��p'�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1����H����lS��h�Oʆ�������8���L�ƨ�D��^����u�<�;�9�#�-�F܁�����^�=��*����
����u�FϺ�����O��N�����4�u�8�
��(�B���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�
�0�
�o�n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h��@���%�u�u����>���<����N��
�����e�n�u�u�$�:����K����lU��N�&���������W��Y����G	�UךU���<�;�9����9�������l��N��1��������}�GϺ�����O��N�����4�u� �������J����	F��s1��2������u�g�9� ���Y����F�D�����6�%�3�
�`��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��^��*���
�m�e�o���;���:����g)��^�����:�e�n�u�w�.����Y����T9��Q��L؊�f�o�����4���:����V��X����n�u�u�&�0�<�W�������A��V�U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Dׁ�����l��N��1��������}�GϺ�����O��N�����4�u�8�
�o�/���O����`2��{!��6�����u�e�3�*����P���F��P ��U���
�d�
� �`�k����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N����l�'�2�f�`�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��a��*ӊ� �b�e�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����C9��[\��*���
�m�c�o���;���:����g)��_����!�u�|�_�w�}����ӗ��9��hY�*��o������!���6�����Y��E��u�u�&�2�6�}��������^��N��1��������}�GϺ�����O��N�����4�u�8�
�e�����A���5��h"��<������}�w�2����I��ƹF��^	��ʧ�<�<�
� �o�k����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���'�2�f�l�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���m�g�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƿ�_9��G\�����f�l�u�u���8���&����|4�Y�����:�e�n�u�w�.����Y����G��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CT��E��F��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l ��^�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	�ӓ�V��^�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�4�-�(���@�ޓ�F��d:��9�������w�m��������l�N�����u�6�%�
�2��N��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
� �l�a�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h[�����f�g�u�u���8���&����|4�N�����u�|�_�u�w�4����+����9��[1�����
�d�3�
�g�e����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��<�����4�9�:�0���F�������F��d:��9�������w�m��������l�N�����u�4�2�d�6�1����&����l ��_�*��o������!���6�����Y��E��u�u�&�2�6�}����H����l	��D1��ۊ�0�
�l�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���:�
�
�d�1��F���	����`2��{!��6�����u�e�3�*����P���F��P ��U���2�d�4�9�-�/����¹��T9��^��U���
���
��	�%���Y����G	�UךU���<�;�9�%�f�m�ށ�����9��T��!�����
����_�������V�=N��U���;�9�%�d�g�4�(���&����\��c*��:���
�����}�������9F������%��9�
��(�F��&���5��h"��<������}�d�9� ���Y����F�D�����
�4�g�a�%�:�D��Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����<�
�&�$���ց�
����	F��s1��2���_�u�u�<�9�1��������W9��N�7�����_�u�w�4��������lW��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������9��E��F���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������G9��P1�C���u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����U��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�o�(���&����\��c*��:���
�����}�������9F�������;�0�
�;�����K����F9��]��F��������4���Y����\��XN�N���u�&�2�4�w�<��������]��1�����f�b�u�u���8���&����|4�N�����u�|�_�u�w�4����+����9��[1�����g�<�3�
�`�d����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��<�����4�9�/�'�$�o�������� F��d:��9�������w�m��������l�N�����u�0�0�0��3����&����l��N��1��������}�GϺ�����O��N�����4�u�0�0�2���������
^��N��1��������}�GϺ�����O��N�����4�u�-�
�2�0�(��&����lT��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�%�(�������9��E��F��u�u��
���(���-���Q��X����n�u�u�&�0�<�W����ԓ�9��h\�L���u�u��
���(���-���U��X����n�u�u�&�0�<�W����ԓ�9��P1�L���u��
����2���+������Y��E��u�u�&�2�6�}��������B9��h��E���8�l�o����0���s���@��V�����2�7�1�g�`�g�5���<����F�D�����8�
�f�
�2��G��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��#���
�e�3�
�d�m����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N��#���
�e�'�2�c�l�W���-����t/��a+��:���g�u�:�;�8�m�L���Yӕ��]��X�����
�
� �g�f��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��X�����
�
�0�
�g�e�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��S�����g�3�
�a�a�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Y
�����
�
�0�
�g�n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��S�����g�;�!�3��i�O���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����3�:�
�
�8�����I���5��h"��<������}�w�2����I��ƹF��^	��ʥ��9�
�d�1��C���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʥ��9�
�d�%�:�C��Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����<�
�&�$����������F��d:��9����_�u�u�>�3�Ͽ�&����Q��]�Oʗ����_�w�}����ӏ��CU��B1�Cފ�g�o�����4���:����V��X����n�u�u�&�0�<�W���	����T9��^��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�e�(���K����CT�=��*����
����u�W������]ǻN�����9�!�%�m��8�(��L����g"��x)��*�����}�u�8�3���B�����Y�����!�%�m�3��k�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�a�
�0��m�E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����e�3�
�c�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R�����
�0�
�e�n�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��G���
�c�g�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���
�e�a�o���;���:����g)��^�����:�e�n�u�w�.����Y����@9��D�����!�'�
�a��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʠ�
�&��&��)��������9��P1�B���u��
����2���+����W	��C��\�ߊu�u�<�;�;�<�(���&����l5��D�*���
�d�o����0���s���@��V�����2�7�1�g�`�g�5���<����F�D�����<�;�<�
��8�(��M����g"��x)��*�����}�u�8�3���B�����Y�����9�
�e�'�0�i�N���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����
�0�
�e�b�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��Z�����m�b�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9�� 1����e�u�u����>���<����N��
�����e�n�u�u�$�:��������9��P1�E���u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���@����lR��N�&���������W������\F��d��Uʦ�2�4�u�8��h�(���&����\��c*��:���
�����}�������9F�������;�0�
�;�����J����_��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�6�:�E�������@9��E��A��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1�%���¹��_9��R��*���g�a�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�`�'�2�c�o�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��V ��D���9�/�'�&�c�;�(��N����	F��s1��2������u�g�9� ���Y����F�D�����4�2�d�4�;�'����M����lR��N�&���������W������\F��d��Uʦ�2�4�u�<�9�4�(݁����� Q�=��*����
����u�W������]ǻN�����9�%��9��o����M����	F��s1��2������u�d�}�������9F������$�<�
�
�2��F��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����a�3�
�l�n�-�W���-����t/��a+��:���g�u�:�;�8�m�L���Yӕ��]��C��D���'�2�a�`�w�}�#���6����e#��x<��G���:�;�:�e�l�}�Wϭ�����G��[�����a�`�u�u���8���&����|4�N�����u�|�_�u�w�4��������P��R	��D��o������!���6�����Y��E��u�u�&�2�6�}����L˹��T9��V��U���
���
��	�%���Y����G	�UךU���<�;�9�%��.����&����W��T��!�����
����_�������V�=N��U���;�9�%��$�1�(ہ�����^�=��*����
����u�W������]ǻN�����9�%��9���F���&����l��N��1��������}�D�������V�=N��U���;�9�%��;��(�������^��N��1��������}�D�������V�=N��U���;�9�4�
�>�����*����U��D��G�������W�W���������D�����f�`�o����9�ԜY�ƿ�T�������`�
� �f�b��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������`�
�0�
�f�m�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��{1��*���0��'�6�"�8�F�������S��N�&���������W��Y����G	�UךU���<�;�9�<��)�4���&����P��R1�D���2�a�l�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƭ�l��h�����
�!�a�3�:�l�W���-����t/��=N��U���;�9�4�
�>�����H����q)��r/�����u�<�;�9�>�����
����A��B��D���3�
�`�a�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��6���
�!� �!�%��@ׁ�����W�=��*����
����u�FϺ�����O��N�����4�u��6��<��������A��V�����3�
�`�a�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������T������'�6� �2�l�O���
����T9��X��U���
���
��	�%���Y����G	�UךU���<�;�9�4��4�(�������@��h��*���o������}���Y����R
��G1�����1�f�l�o���2���s���@��V�����3�
�`�b�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������1����d�u�u����>���<����N��S�����|�_�u�u�>�3�Ϸ�&����\��X��D���3�
�c�m�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������[�����:�%�d�c�%�:�C��Y�Ɵ�w9��p'��#����u�d�1� �)�W���s���@��V�����2�6�0�
��.�F؁�
����\��c*��:���n�u�u�&�0�<�W���
����W��_��U�����n�u�w�.����Y����V��Q��C���%�u�u����>���<����N��
�����e�n�u�u�$�:��������9��P1�G���u��
����2���+������Y��E��u�u�&�2�6�}��������F9��\��G��������4���Y����\��XN�N���u�&�2�4�w�)�G��L����l��N��1��������}�D�������V�=N��U���;�9�9�
��i�(���&����l��hZ�C��������4���Y����W	��C��\�ߊu�u�<�;�;�<�(���&����l5��D�*���
�m�o����0���s���@��V�����2�7�1�f�b�g�5���<����F�D�����!�e�a�`�2�l����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*������0�:�o�E���H����lR��N�&���������W��Y����G	�UךU���<�;�9�7�1�m�F��&����V��T��!�����
����_�������V�=N��U���;�9�7�3�g�l�Cց�����`2��{!��6�ߊu�u�<�;�;�?����H����BV�=��*����
����u�FϺ�����O��N�����4�u� �
��o�N�������F��d:��9�������w�l��������l�N�����u� �
�
�e�d���Cӵ��l*��~-�U���&�2�4�u�"��(��@����\��c*��:���n�u�u�&�0�<�W���&ù��_��N�&���������W��Y����G	�UךU���<�;�9�9���Cځ�&ù��W��D^��U���
���
��	�%���Y����G	�UךU���<�;�9�9���Cځ�&ù��F��d:��9����_�u�u�>�3�ϲ�&ù��9��1�����&�u�u����>���<����N��S�����|�_�u�u�>�3�ϲ�&ù��9��1��D�������W�W�������
��1�@���e�"�d�o���;���:���F��P ��U���e�a�`�0�g�9�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��[��*��
�
�
�d�m��3���>����v%��eN��Eʱ�"�!�u�|�]�}�W�������G9��Z�����4�1�0�&�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������G9��Z�����6�e�o����0���s���@��V�����a�`�0�d�6�9����Y�Ɵ�w9��p'��#����u�d�1� �)�W���s���@��V�����a�`�0�d�4�l�Mύ�=����z%��N�����4�u�!�e�c�h�������5��h"��<��u�u�&�2�6�}����M�ӓ�lW��N�&���������W��Y����G	�UךU���<�;�9�9���Cځ�&¹��\��c*��:���
�����l��������l�N�����u��9�
�8�����
����lR��T��!�����
����_�������V�=N��U���;�9�4�
�>�����*����^��D��B�������W�W���������D�����a�g�o����9�ԜY�ƿ�T�������6�0�
��$�l�(���&���5��h"��<��u�u�&�2�6�}��������lR��T��:����n�u�u�$�:����	����l��F1��*���e�3�8�d�w�}�#���6����9F������4�
�<�
�3��C���Y����v'��=N��U���;�9�<�
�#���������F��V�����`�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��1��*��m�%�u�u���8���&����|4�^�����:�e�n�u�w�.����Y����@��h��A���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l ��W�����u��
����2���+������Y��E��u�u�&�2�6�}��������U��\��A��������4���Y����W	��C��\�ߊu�u�<�;�;�)��������9��T��!�����
����_������\F��d��Uʦ�2�4�u�8�����I����	F��s1��2������u�a�}�������9F������!�%�m�
�6�)����&����R��N�&���������W��Y����G	�UךU���<�;�9�0�'�����KŹ��\��c*��:���
�����l��������l�N�����u�8�
�d�1��A݁�K����g"��x)��*�����}�d�3�*����P���F��P ��U���
�g�3�
�a��C��*����|!��h8��!���}�e�1�"�#�}�^�ԜY�ƿ�T��
�����;�d�3�
�o��F��*����|!��h8��!���}�f�1�"�#�}�^�ԜY�ƿ�T�������d�3�
�m��l�Mύ�=����z%��r-��'���f�1�"�!�w�t�}���Y����R
��O�����
�
� �c�g�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��C��F܊� �c�e�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����G��_�����g�
�d�o���;���:����g)��[����!�u�|�_�w�}����Ӓ��lU��Q��Gފ�f�o�����4���:����S��S�����|�_�u�u�>�3�Ϯ�+����G9��Q��F؊�d�o�����4���:����S��S�����|�_�u�u�>�3�ϳ�����l ��]�����u��
����2���+������Y��E��u�u�&�2�6�}����Hǹ��lS��h�Oʆ�������8���O�ƨ�D��^����u�<�;�9���(���O�Г�F��d:��9�������w�l�W������]ǻN�����9���
���(���O�ԓ�F��d:��9�������w�m��������l�N�����u�8�
�l�1��Aׁ�K����g"��x)��*�����}�d�3�*����P���F��P ��U���
�e�3�
�`��E��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������d�3�
�m��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��V ��*܊� �c�g�%�w�}�#���6����e#��x<��@���:�;�:�e�l�}�Wϭ�����@��Z��*���!�3�
�m��l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��Z��@���
�d�
�d�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������^��1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������Q��B1�M���u�u��
���(���-���Q��X����n�u�u�&�0�<�W���&�ѓ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��o����I����\��c*��:���
�����}�������9F������!�%�d�m�1��Eہ�H����g"��x)��*�����}�b�3�*����P���F��P ��U���
� �b�m�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�*���b�a�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h�����
�b�
�d�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������^��1��*���
�g�o����0���/����aF�
�����e�n�u�u�$�:��������9��hY�*��o������!���6�����Y��E��u�u�&�2�6�}����M����_��G\��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�:��Eށ�����l��N��1��������}�BϺ�����O��N�����4�u�8�
�b�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʥ�:�d�3�
�f��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��D���3�
�d�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��\�����g�
�d�o���;���:����g)��[����!�u�|�_�w�}����Ӓ��lW��h��M���%�u�u����>���<����N��
�����e�n�u�u�$�:����&����_��h��M���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l �� W�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����T��N�&���������W������\F��d��Uʦ�2�4�u�8��o�(���A�ԓ�F��d:��9�������w�m��������l�N�����u�
�
� �o�e����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���3�
�l�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��M���
�m�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��1��*��
�a�o����0���/����aF�
�����e�n�u�u�$�:��������U��\��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_�������V�=N��U���;�9�!�%�o���������U��Z��F��������4���Y����W	��C��\�ߊu�u�<�;�;�8����H����W��G\��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�:��O���&����CT�=��*����
����u�FϺ�����O��N�����4�u�8�
�d����A����	F��s1��2������u�f�}�������9F������%�&�
�
�"�d�C���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����
�
� �l�c�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��C��D���3�
�b�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����C	��h_�����3�
�`�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������hX�����m�
�d�o���;���:����g)��[����!�u�|�_�w�}����Ӓ��lP��Q��MҊ�g�o�����4���:����S��S�����|�_�u�u�>�3�ϲ�&¹��l_��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2�o����N˹��\��c*��:���
�����}�������9F������!�%�
� �n�e����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*��
� �d�d��n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���d�g�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƾ�EU��B1�DҊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���K�ד�R��Q��Cڊ�d�o�����4���:����U��S�����|�_�u�u�>�3�Ϫ�	����U��]�����u��
����2���+������Y��E��u�u�&�2�6�}����K����l ��^�*��o������!���6��� F��@ ��U���_�u�u�<�9�1����H����V��h�Oʆ�������8���L�ƨ�D��^����u�<�;�9�8�����Hƹ��l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}����K����l	��D1�����e�g�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӵ��T��V�����
�
� �d�g��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��C݊� �d�b�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����a��R_�����0�:�
�
�"�l�Oہ�K����g"��x)��*�����}�u�8�3���B�����Y��'���0�
�9�
�2�2�(܁�����9��T��!�����
����_�������V�=N��U���;�9�!�%�a���������9��T��!�����
����_�������V�=N��U���;�9�!�%�a����@Ź��\��c*��:���
�����}�������9F������&�9�!�%�a�;�(��I����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�f��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʺ�
�:�1�d��l����I�Г�F��d:��9�������w�m��������l�N�����u�4�2�d�6�1����&����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����A����W��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��l�(�������^��N�&���������W������\F��d��Uʦ�2�4�u�
�e��F���&����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�n�(���H����CU�=��*����
����u�W������]ǻN�����9�!�%�d�b�;�(��M����	F��s1��2������u�g�9� ���Y����F�D�����8�
� �d�`��D��*����|!��h8��!���}�g�1�"�#�}�^�ԜY�ƿ�T�������!�c�3�
�f�h����Y����)��t1��6���u�`�u�:�9�2�G��Y����Z��[N�����d�3�
�d�n�-�W���-����t/��a+��:���`�u�:�;�8�m�L���Yӕ��]��C��F���
�g�g�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����G��1��*��b�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����^��B1�D؊�f�o�����4���:����W��S�����|�_�u�u�>�3�ϳ�����F9��[��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.�(���&����l ��\�*��o������!���6���F��@ ��U���_�u�u�<�9�1����K����T��h�Oʆ�������8���L�ƨ�D��^����u�<�;�9�#�-�C���&����l��N��1��������}�B�������V�=N��U���;�9�!�%�f����K˹��\��c*��:���
�����n��������l�N�����u�8�
�e�1��E���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʡ�%�d�
� �f�k�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
� �d�f��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���d�`�
�d�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������lT��1��*��m�%�u�u���8���&����|4�]�����:�e�n�u�w�.����Y����R��B1�Lي�g�o�����4���:����W��S�����|�_�u�u�>�3�Ϫ�	����P��h��D��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������9��h_�B���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����K˹��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Fف�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��i����J�Փ�F��d:��9�������w�h��������l�N�����u�8�
�b�1��D���	����`2��{!��6�����u�e�3�*����P���F��P ��U���%�3�
�f�`�-�W���-����t/��a+��:���`�1�"�!�w�t�}���Y����R
��Z��F���
�f�f�%�w�}�#���6����e#��x<��@ʱ�"�!�u�|�]�}�W�������^��1��*��d�%�u�u���8���&����|4�]�����:�e�n�u�w�.����Y����W��B1�@ߊ�g�o�����4���:����S��S�����|�_�u�u�>�3�Ϯ�+����G9��Q��F���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l ��]�*��o������!���6�����Y��E��u�u�&�2�6�}����A����U��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��<�E�������_��N�&���������W��Y����G	�UךU���<�;�9�!�'�k�(���H����CW�=��*����
����u�W������]ǻN�����9�'�3�
�d�n����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*��� �d�l�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����B��B1�Dڊ�f�o�����4���:����V��X����n�u�u�&�0�<�W�������]9��Q��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����U��^�����u��
����2���+������Y��E��u�u�&�2�6�}�(���K�Փ�F9��Y��G��������4���Y����W	��C��\�ߊu�u�<�;�;�)��������U��N�&���������W������\F��d��Uʦ�2�4�u�0��0�O���&����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�d����M�ӓ�F��d:��9�������w�m��������l�N�����u�8�
�d�1��D���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�`�3��i�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�b�3�
�c�l����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N�����%�d�3�
�c�i����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���d�
� �d�a��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����e�3�
�a�a�-�W���-����t/��a+��:���g�u�:�;�8�m�L���Yӕ��]��D�����a�3�
�a�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��*���d�f�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G_�����a�l�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lT��Q��G���%�u�u����>���<����N��
�����e�n�u�u�$�:��������CW��Q��A���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l ��Z�*��o������!���6�����Y��E��u�u�&�2�6�}���H����\��Y1��*��f�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������U��W�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�-�ށ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�:�e�;�(��I����	F��s1��2������u�f�}�������9F������!�%�m�
�"�l�C܁�J����g"��x)��*�����}�u�8�3���B�����Y�����
�4�!�3��h�A���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����g�
� �d�b��F��*����|!��h8��!���}�f�1�"�#�}�^�ԜY�ƿ�T����*���3�
�`�d�'�}�W���&����p9��t:��U���u�:�;�:�g�f�W���
����_F��h��D��
�d�o����0���/����aF�
�����e�n�u�u�$�:��������lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�(���H����CT�=��*����
����u�W������]ǻN�����9�!�%�d�g�;�(��J����	F��s1��2������u�g�9� ���Y����F�D�����8�
�b�3��h�@���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����3�
�`�d�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������1����� �d�g�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h\�����c�l�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƞ�]��h8��*���d�d�
�g�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������l0��B1�Dӊ�g�o�����4���:����S��S�����|�_�u�u�>�3�ϱ�&����W��^1��*��f�%�u�u���8���&����|4�N�����u�|�_�u�w�4����+����9��[1����� �d�g�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����a��R\�����;�&�d�<�1��A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���2�d�4�9�8�8�(ށ�����9��T��!�����
����_�������V�=N��U���;�9�!�%�d����L¹��\��c*��:���
�����}�������9F�������;�0�
�;�����&����S��G\��U���
���
��	�%���Y����G	�UךU���<�;�9��9�8�(���&����@9��Q��C���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����]	��Q��C���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����U��X�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	�Г�F9��]��G��������4���Y����\��XN�N���u�&�2�4�w�8�(���HĹ��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�8�����HĹ��U��]�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�����&����\��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CW��Q��B���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϯ�H�ߓ�l ��X�*��o������!���6�����Y��E��u�u�&�2�6�}�(��&����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����@����Q��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����U�� ]�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)�܁����� 9��T��!�����
����_�������V�=N��U���;�9�6�'�.�l��������Q��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�6�:�E�������@9��Y�����
�b�`�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��_�� ��b�
�f�o���;���:����g)��^�����:�e�n�u�w�.����Y����A��]��*���d�c�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�g�8�-�>�;�(��N����	F��s1��2������u�g�9� ���Y����F�D�����
�g�
�
�"�l�Oށ�K����g"��x)��*�����}�u�8�3���B�����Y�����&�<�;�f�1��@���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�b�3�
�`�d����Y����)��t1��6���u�d�u�:�9�2�G��Y����Z��[N��#���
�
� �d�g��E��*����|!��h8��!���}�b�1�"�#�}�^�ԜY�ƿ�T����*���f�
� �d�f��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����g�3�
�m�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����
� �d�f��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�m�e�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��[1�����3�
�m�b�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�M���
�m�m�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��1�����4�
� �d�b��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��*���d�`�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƽ�e��h_�����m�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ư�A��1��*���d�c�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��GW�����3�
�m�g�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������1��*��m�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������lW��X��D���
�m�f�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������R��1�����0�
�
�:��l����A�ߓ�F��d:��9�������w�m��������l�N�����u�'�0�2�f�n�ށ�����9��T��!�����
����_�������V�=N��U���;�9��;�2���������l��h�����l�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӵ��T��V�����
�
�d�d��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʱ�9�!�1�:�2��(���H����CU�=��*����
����u�W������]ǻN�����9�&�9�!�'�m����@�Փ�F��d:��9�������w�m��������l�N�����u�0�&�2�5�)�F���&����l��N��1��������}�GϺ�����O��N�����4�u�8�d��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʦ�9�!�%�g�1��N���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�l�3�
�n�j����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���a�
� �d�b��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��S�����/�'�&�d�1��O���	����`2��{!��6�����u�e�3�*����P���F��P ��U���0�0�
�0�8��(���&����
P��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�1�;�)��������l��h�����l�f�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӄ��V��h�����l�m�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lQ��Q��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϻ�����l	��D1��ۊ� �d�f�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����Q��E	��Gۊ�0�:�2�;�>����@ƹ��\��c*��:���
�����}�������9F������&�2�
�&�>�3�F���&����l��N��1��������}�GϺ�����O��N�����4�u�'�0�0�l�F���&����V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9� �3�/����H����V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�!�/����H����_��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�>�3��������]	��Q��E���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	�ד�F9��[��G��������4���Y����\��XN�N���u�&�2�4�w�/����&����l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}����I����V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��<�E�������S��N�&���������W��Y����G	�UךU���<�;�9�&�;�)���&����A��h��G��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CR��Q��E���%�u�u����>���<����N��
�����e�n�u�u�$�:��������VW��B1�Fۊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����9��h\�B���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����K����V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����^��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�%��1�(�������F9��Y��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.����	�ғ�F9��W��F��������4���Y����W	��C��\�ߊu�u�<�;�;�����&����\��h\��*���3�
�d�c�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��Gڊ� �g�d�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��h��G��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CT��Q��D���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����U��_�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	�ד�F9��_��G��������4���Y����\��XN�N���u�&�2�4�w�8����&����@9��h\�D���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������V��h ��*���g�a�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƨ�_��S1�����e�;�!�<�1��F���	����`2��{!��6�����u�e�3�*����P���F��P ��U���0�2�
�
�"�o�Bց�K����g"��x)��*�����}�u�8�3���B�����Y�����f�
� �g�a��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��S�����:�0�
�
��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʷ�8�'�0�g��8��������F9�� [��G��������4���Y����\��XN�N���u�&�2�4�w�4����
����U��Z�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�?��������Z9��h\�E���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l ��_�*��o������!���6�����Y��E��u�u�&�2�6�}��������F9��W��G��������4���Y����\��XN�N���u�&�2�4�w�4����
����]	��Q��D���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	ƹ��lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�5�0��������F9��\��G��������4���Y����\��XN�N���u�&�2�4�w�0�(������� V��N�&���������W������\F��d��Uʦ�2�4�u�
�6�o�B���&����l��N��1��������}�E�������V�=N��U���;�9�&�9�#�-�N�������]9��h\�G���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l ��\�*��o������!���6��� F��@ ��U���_�u�u�<�9�1��������F9��^��G��������4���Y����\��XN�N���u�&�2�4�w�8�(���Kƹ��lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�(���K����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�k����K�ғ�F��d:��9�������w�m��������l�N�����u�
�4�g�b�0����&����l��N��1��������}�E�������V�=N��U���;�9�&�9�#�-�C���&����l��N��1��������}�E�������V�=N��U���;�9�%��;��@���&����l��N��1��������}�D�������V�=N��U���;�9�!�%�f�d����J�ד�F��d:��9�������w�e��������l�N�����u�8�
�a��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʧ�g�3�
�f�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h��G���
�f�a�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������Q��Q��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϯ�&����T��h��G��
�g�o����0���/����aF�
�����e�n�u�u�$�:����&����lT��Q��G���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l ��]�*��o������!���6��� F��@ ��U���_�u�u�<�9�1��������G9��Q��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����l ��]�*��o������!���6�����Y��E��u�u�&�2�6�}����L����U��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��8����Hǹ��G9��h\�C���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������F9��V��F��������4���Y����\��XN�N���u�&�2�4�w�2�(�������lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�4�/����&����l��N��1��������}�GϺ�����O��N�����4�u�0�0�2�����&����lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'�3��������P��N�&���������W������\F��d��Uʦ�2�4�u�'�2�:�(�������T��N�&���������W������\F��d��Uʦ�2�4�u�8��k����J�ғ�F��d:��9�������w�m��������l�N�����u�
�m�<�1��C���	����`2��{!��6�����u�e�3�*����P���F��P ��U���0�2�a�
�2�2��������R��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:�o�B�������]9��h\�E���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����J����R��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��D���&����l��N��1��������}�GϺ�����O��N�����4�u�-�
��%��������G��V��*���&�3�
�a�c�-�W���-����t/��a+��:���g�u�:�;�8�m�L���Yӕ��]��U�����<�<�
� �e�j�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��#���
�f�8�-�1��C���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʥ��9�
�
�"�o�O؁�J����g"��x)��*�����}�f�3�*����P���F��P ��U���
�a�
� �e�m�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
� �g�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1��&���!��&�9�#�����&�ߓ�l ��[�*��o������!���6��� F��@ ��U���_�u�u�<�9�1����8����F��U�� ����9�0�l�����Oʹ��\��c*��:���
�����n��������l�N�����u�-�
��/�(�(�������l0��B��L���3�
�`�c�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��C1��*���a�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������K!��x��2���!�'��
�&�<�(�������9��T��!�����
����_�������V�=N��U���;�9�7�:���G���&����G��x�����
�
� �g�g��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��U��*���e� �
�'�6�8�(���<����l��B1�@ފ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����U��[�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����R��GZ��U���
���
��	�%���Y����G	�UךU���<�;�9�'�!����Nù��\��c*��:���
�����}�������9F������&�9�!�%�`�;�(��M����	F��s1��2������u�g�9� ���Y����F�D�����6�%�b�;�#�;�(��K����	F��s1��2������u�g�9� ���Y����F�D�����8�
�l�3��h�A���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�a�
� �e�l�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�`�
�0�8�:����&����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�l�O�������]9��h\�E���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Aù��lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����H����P��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�/���������R��a1��*��m�%�u�u���8���&����|4�Z�����:�e�n�u�w�.����Y����]	��h�����c��3�
�a�j����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N�����1�
�0�8�b�l�!���&����l��N��1��������}�E�������V�=N��U���;�9�:�
�8�9����O�Փ�F��d:��9�������w�m��������l�N�����u�0��9�1��A���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʺ�
�:�1�
�"�o�Oہ�K����g"��x)��*�����}�u�8�3���B�����Y�����:�1�
� �e�d�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����d�3�
�c�o�-�W���-����t/��a+��:���g�u�:�;�8�m�L���Yӕ��]��Q�����
�0�8�a�`�����O�ד�F��d:��9�������w�o�W������]ǻN�����9�;�"�0�d�;�(��I����	F��s1��2������u�e�}�������9F������;�"�0�`�1��@���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʻ�"�0�a�3��j�@���Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����0�l�3�
�`�e����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N�����f�a�6�&��(�E��&���5��h"��<������}�c�9� ���Y����F�D�����0��9�
�"�o�Aہ�J����g"��x)��*�����}�a�3�*����P���F��P ��U����9�
� �e�h�(��Cӵ��l*��~-��0����}�a�1� �)�W���s���@��V�����8�`�
� �e�e�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
�c�c�%�w�}�#���6����e#��x<��Gʱ�"�!�u�|�]�}�W�������V
��Z�*���g�l�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G[�����b�b�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӗ��R
��1��*��g�%�u�u���8���&����|4�Z�����:�e�n�u�w�.����Y����_T��h��G��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������9��h\�A���u�u��
���(���-���S��X����n�u�u�&�0�<�W���&�Փ�F9��^��D��������4���Y����W	��C��\�ߊu�u�<�;�;�-�!���&ƹ��l ��Y�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������l ��Y�*��o������!���6���F��@ ��U���_�u�u�<�9�1����AŹ��lT��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������R��N�&���������W��Y����G	�UךU���<�;�9�'��i����A�ޓ�F��d:��9�������w�o�W������]ǻN�����9�3�%�-��	�8���4����C
��\��#���
�m�`�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����G��V�� ��a�
�d�o���;���:����g)��[����!�u�|�_�w�}����Ӏ��l��{:�� ��� �!�%�,�f�i�!���&����l��N��1��������}�E�������V�=N��U���;�9�'��b�;�(��K����	F��s1��2������u�e�}�������9F������3�%�-� ����������J9�� 1�����m�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�C9��b"��:����9�<�9��o�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�-���;�������_��[��Gފ�
� �g�a��o�Mύ�=����z%��r-��'���c�1�"�!�w�t�}���Y����R
��h<�� ���&�d�
� �e�l�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��'���9�
�
� �e�n�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����� ���!��1����&����e9��h\�@���u�u��
���(���-���P��X����n�u�u�&�0�<�W���&����T��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�'�>�4�(���J����CT�=��*����
����u�W������]ǻN�����9�$�
�&�>�3�@���&����l��N��1��������}�GϺ�����O��N�����4�u�8�
�g�;�(��K����	F��s1��2������u�d�}�������9F������%��9�
�f�;�(��O����	F��s1��2������u�d�}�������9F������;�"�<�;�>��(���J����CU�=��*����
����u�W������]ǻN�����9�!�%�l��(�D��&���5��h"��<������}�w�2����I��ƹF��^	��ʶ�'�,�d�3��m�B���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����g�3�
�e�a�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��hZ��ۊ� �f�m�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����W��C�����&�f�3�
�g�m����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������d�3�
�e�o�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E�����f�3�
�d�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��F���
�d�e�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��R
�����g�3�
�e�a�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h]��ۊ� �f�l�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����Q��E	��E���8�'�4�
�f�;�(��H����	F��s1��2������u�g�9� ���Y����F�D�����8�g�b�1�:�/��������9��T��!�����
����_�������V�=N��U���;�9�!�%�c�;�(��J����	F��s1��2������u�g�9� ���Y����F�D�����;�0�3�:�����Jʹ��\��c*��:���
�����}�������9F������:�0�3�:�����Hƹ��\��c*��:���
�����}�������9F������!�%�`�3��l�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����2�
�
�f�1��F���	����`2��{!��6�����u�e�3�*����P���F��P ��U���0�3�:�
��2�(���J����CT�=��*����
����u�W������]ǻN�����9�%��9��m�(���&����P��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u��<�E���Kù��lU��1��U����
�����#���Q����\��XN�N���u�&�2�4�w��(���J����CT�=��*����
����u�W������]ǻN�����9�'�<�<��(�D��&���5��h"��<������}�w�2����I��ƹF��^	��ʤ�
�&�<�;�n�;�(��O����	F��s1��2������u�g�9� ���Y����F�D�����8�
�a�3��o�F���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����9�
�f�3��o�B���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����<�;�<�
��(�D��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�l�
� �d�l�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����g�3�
�g�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��V ��D���9�:�0�
��(�D��&���5��h"��<������}�w�2����I��ƹF��^	��ʇ�;�0�
�9��8����&����U��G\��U���
���
��	�%���Y����G	�UךU���<�;�9��9�8�(���&����lR��B1�Gӊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&�Г�F9��\��G��������4���Y����\��XN�N���u�&�2�4�w��F���&����S��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�1�;�)��������l ��\�*��o������!���6�����Y��E��u�u�&�2�6�}�(���&�ԓ�F9�� Y��G��������4���Y����\��XN�N���u�&�2�4�w�/����&�ғ�F9��]��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������_��N�&���������W������\F��d��Uʦ�2�4�u�0�2�8�(���
�Փ�F9��]��F��������4���Y����\��XN�N���u�&�2�4�w��O���&����Q��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�7�:�/��������T��^\�� ��e�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����
_��R�����3�
�f�c�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������X�� ��d�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����A ��@1�����f�m�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӊ��A ��@1�����g�a�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��Q��B1�Gӊ�g�o�����4���:����V��X����n�u�u�&�0�<�W�������Z9��h��F��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������_	��1�����
�f�`�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������l0��1�@���-�3�
�f�f�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��G1��؊�
�g�3�
�d�d����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����3�
�f�`�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h �����'�
�f�
�"�n�Aց�K����g"��x)��*�����}�d�3�*����P���F��P ��U���
�m�3�
�d�i����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*����&�
�!�"�)����N˹��U��V�����u��
����2���+������Y��E��u�u�&�2�6�}�;���&����l5��B�����b�
�
� �d�e�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����l�3�
�f�o�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��Eڊ� �f�e�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��C���
�a�m�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�L���8�'�4�
�"�n�D߁�K����g"��x)��*�����}�u�8�3���B�����Y�����d�d�3�
�c�e����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���`�
� �f�d��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����a�
�0�:�0�3����M�ޓ�F��d:��9�������w�m��������l�N�����u�8�
�e��(�D��&���5��h"��<������}�w�2����I��ƹF��^	��ʦ�9�!�%�e�1��C���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�c�
�"�n�A߁�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�l�3��i�E���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�`�
� �d�o�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*����&�
�!�"�)����Aƹ��U��W�����u��
����2���+������Y��E��u�u�&�2�6�}�����Փ�F9�� Z��G��������4���Y����\��XN�N���u�&�2�4�w�8�$���&����P��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�2��ׁ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�'�4�3�C���&����l��N��1��������}�GϺ�����O��N�����4�u�'�6�9�h����L�ߓ�F��d:��9�������w�m��������l�N�����u�0��9�f�;�(��H����	F��s1��2������u�d�}�������9F������;�"�0�d��(�D��&���5��h"��<������}�f�9� ���Y����F�D�����0��9�g�1��B���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʻ�"�0�d�
�"�n�Dށ�J����g"��x)��*�����}�d�3�*����P���F��P ��U����9�`�3��h�A���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����0�d�
� �d�n�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����9�c�3�
�b�o����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����d�
� �f�`��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�� ��&���b�3�
�`�g�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��C��D���3�
�c�m�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h_�*���f�a�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��1��*��l�%�u�u���8���&����|4�^�����:�e�n�u�w�.����Y����l
��q��9���
�
� �f�b��D��*����|!��h8��!���}�e�1�"�#�}�^�ԜY�ƿ�T����*��
� �f�g��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����
�c�l�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������l��[�����:�%�6�&��(�D��&���5��h"��<������}�f�9� ���Y����F�D�����
�
��9��2�(���	����F9��\��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.����	����lU��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����&����^��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)�ށ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�0�n�;�(��O����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�c�1��@���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�a�3��k�D���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����0�8�
�;��3��������A��1��*��`�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����`3��x��G���3�
�b�f�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��9����!�g�g�1��@���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ��9�
�b�1��@���	����`2��{!��6�����u�d�w�2����I��ƹF��^	��ʲ�%�3�
�b��8�Mύ�=����z%��N�����4�u�%�&�0�>����-����l ��h_��U���
���n�w�}�����ƭ�l��h��*��c�o�����}���Y����R
��G1�����0�
��&�d�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������F��u!��0���_�u�u�<�9�1��������V��c1��A���8�f�o����0���s���@��V�����2�7�1�g�d�}�W���5����9F������4�
�<�
�$�,�$���ƹ��^9��N��1�����_�u�w�4��������T9��S1�F���u����l�}�Wϭ�����R��^	������
�!�
�$��W���-����t/��=N��U���;�9�4�
�>�����H���$��{+��N���u�&�2�4�w�/�(���M�Г�VF��d:��9����_�u�u�>�3�Ͽ�&����@�=��*����
����u�NϺ�����O��N�����4�u�%�&�0�?���Y�Ǝ�|*��yUךU���<�;�9�4��4�(���&���$��{+��N���u�&�2�4�w�-��������F��u!��0���_�u�u�<�9�1��������W9��T��:����n�_�u�w�2�����ơ�"�� V��*ڊ�1�#�f�;��o���&�ƅ�9F�	�����u�_�u�u�w�}�3��0����v4��N��U��������g�>���>����F�N�����
���u�w��2���B���F�
��D�����o����%�ԜY���F��B��<���u�u����}�L���YӖ��GF�N��U���6�>�o��w�	�(���0��ƹF�N�����u�u�����0���s���F�S��U���������!���6���F��@ ��U���_�u�u�u�w�4�F��0�Ɵ�w9��p'��#����u�f�u�8�3���B���F���Oʜ�u��
���f�W���Y����\��N��!ʆ�������8���J�ƨ�D��^��\�ߊu�u�;�u�8�-����B��ƹF��X�����u���d�o�;�G���������Z��U���u�u�2�;�%�>�_���Y���/��N��!����_�u�u�w�}�"���-����	F��c+��'�ߊu�u�u�u�>�m� ���1����}2��r<�U���u�u�1� ���#���Y����t#��UךU���:�!�}�u�w�}�WϺ�����z(��c*��:���
�����l��������l�N��Uʱ� �u�u� �w�	�(���0����p2��F�U���;�:�e�u�l�}�Wϻ�Ӆ��C	��Y����u�6�8�:�2�)����<����U9��Z�����d�;�
�m��h�Fϗ�s���T��E��]���u�u�u��w�}�9���<��ƹF�N�� �����u�u���2��Y���F��^ ��"����o�����}���Y���W��h9��!���u����l�}�W���Yӂ��G9��s:��Oʜ����|�]�}�W�����ƹF�N����o��u����>���<����N��
�����e�n�u�u�w�}����Y�ƅ�5��h"��<������}�`�9� ���Y����F�N�����u�u� �u���8���&����|4�Z�����:�e�u�n�w�}��������]��dװU���6�8�:�0�#�0�A���N�Ѫ�9��Q1��D��u��u�u�0�3����Q���F�*�����!�u�u����L���Y���'��E��'���0�o�����}���Y���r��R�����u�u����}�L���YӖ��GF�N��U���6�>�o��w�	�(���0��ƹF�N�����u�u�����0���s���F�V
�����u�u�����0���/����aF�
�����e�n�u�u�w�}���Cӯ��`2��{!��6�ߊu�u�u�u�g�g�8���*����|!��h8��!���}�d�1�"�#�}�^�ԜY���F��S�����u������4���:����W��X����n�u�u�u�w�>�F��0�Ɵ�w9��p'�����u�u�u�0�w�}�9ύ�=����z%��N��U���1�u�u����;���:����g)��]����!�u�|�|�]�}�W���Y����\��CUװ���u�:�%�;�9�}�1ٚ�H����lV��C1��A���0�e��_�w�}�������F�N��1����1�=�o��	�0���s���F�v
�����4�2�u�u���2��Y���F��S
�����1�=�o����%���s���C	��FךU���u�u�9�u�w��$���5����l�N��Uʧ�&�!�o��w�	�(���0��ƹF�N�����&�e�o��w�	�(���0����p2��F����!�u�|�_�w�}�W�������z(��c*��:���n�u�u�u�w�,�W���,�Ɵ�w9��p'��#����u�f�u�8�3���B���F������d�o��u���8���&����|4�N�����u�|�_�u�w�}�W���Y�ƅ�5��h"��<��u�u�u�u� �l�Mϗ�Y����)��tUךU���u�u�d�o��}�#���6����e#��x<��F���:�;�:�e�l�}�W���Yӗ��	F��cN��1��������}�D�������V�UךU���;�u�:�%�9�3�L�ԶY����\��Y��U����d�m�3�g�1�(߁�Mƹ��F��=N��U���0�<�u�_�w�}�W�������W��N��!����_�u�u�w�}����
����T�'��0���n�u�u�u�w�����
����[F��~ ��2���|�_�u�u�8�)�_���Y�����T��;ʆ�����]�}�W���Y����GF��~ ��!�����n�u�w�}�WϿ�����F��~ ��!�����
����_�������V�=N��U���u�0�u�u���3���>����F�N�����u� �u����>���<����N��
�����e�n�u�u�w�}��������	F��=��*����
����u�W������]ǻN��U���0�u�u����;���:���F�N��D���u��
���L���Y�����N��U���
���
��	�%���Hӂ��]��G�U���u�u�$�u�w��W���&����p9��t:��U��u�:�;�:�g�}�L���YӃ����G����_�_�0�<�]�}�W���&ù��_��T�����;�;�u���l�Oظ�I����lV��Z�U���2�;�'�6�:�-�_���Y���"��V9�����k�f�y�u�w�}�Wϟ�����a��RN��U���u�u�u�u��9��������X�d��Uʥ�'�u�4�u�]�}�W���Y����X��G1���ߊu�u�u�u�2�8�W�������GJǻN��U���1�'�&�e�j�}����&����l��E��E�ߊu�u�u�u�2�}�Iϼ��֓�R��T����u�u�u�e�j�}����&����l��=N��U���u�1�'�&�f�`�W���&ù��_��S
����_�u�u�u�w�8�W�������lW��1��D�ߊu�u�u�u�2�}�Iϼ��֓�R��@����u�u�u�d�j�}����&����l��dךU���!�e�a�`�2�m�"������]����1��m�3�e�9���Cځ�&���F��Y��ʸ�%�}�u�u�w�}�3���.����[�_�U���u�u��1�2�.����Y���l�N��Uʔ�1�0�&�<�#�}�I��s���C	����U�ߊu�u�u�u�;�}�IϿ�&����9F�N��U���0�u�k�4��.�[���Y�����E��E��u�!�e�a�b�8�G�������JǻN��U���0�u�k�9���Cځ�&ù��JǻN��U���e�h�u�!�g�i�B���I����9F�N��U���'�&�d�h�w�)�G��L����l��E��D�ߊu�u�u�u�2�}�Iϲ�&ù��9��1��D�ߊu�u�u�u�2�}�Iϲ�&ù��9��1��D�ߊu�u�u�u�f�`�W���I����l��h
����u�u�u�d�j�}����M�ӓ�lV��G����u�!�e�a�b�8�F���CӅ��C	��Y��3ܑ�d�m�3�e�;��(��&����F�P�����8�%�}�u�w�}�WϚ�����G�	N�Y���u�u�u��3�8�������U�N��U����1�0�&�>�)�W���K���F��E�����_�u�u�u�w�1�W�������XJǻN��U���0�0�u�k�6����Y���F��S
����h�u�!�e�c�h��������@��=N��U���u�0�u�k�;��(��&����P��=N��U���u�e�h�u�#�m�C����ד�JǻN��U���1�'�&�d�j�}����M�ӓ�lW��S
����_�u�u�u�w�8�W�������R��R1����_�u�u�u�w�8�W�������R��R1����_�u�u�u�w�l�J����֓�S��h_��D�ߊu�u�u�u�f�`�W���I����l��h�N�ߊu�u�
�
�3�+�Dݰ�&�Ԣ�lU�� 1��U���:�%�;�;�w��3��AĀ��l ��A1����g�&�f�
�]�}�W�������^��d��U���u��u�k�f�W�W���Y�Ƃ�~9��v)��H���y�u�u�u�w�9�߁�0����X�BךU���u�u�<�d� ��?��Y����F�N�����
���u�i�n�^���YӖ��GF��GN��U���u�u�6�>�j�}�������F�N�����h�u�%�'�#�W�W���Y�ƨ�]V�	N��E���
�<�y�u�w�}�WϺ������h�����_�u�u�u�w�8�J�������lR��h�����u�u�u�:�#�`�W���&����V��G����u�
�
�1�!�n����K����9��b_��U���%�;�;�u���F���֓�W��\��*���&�f�
�_�w�}�����ơ�CF�N��U����u�k�d�]�}�W���Y����`2��rN��U���u�u�u�u�3�3�(���-���U��=N��U���u�<�d����J���K���F�N�� �����u�k�d�t�W���	����^��d��U���u�6�>�h�w�-����s���F�E����u�%�'�!�]�}�W���Y����[�G1�����<�y�u�u�w�}����Y����lW��Y1���ߊu�u�u�u�2�`�W���&����P��RBךU���u�u�:�!�j�}��������l��dךU���
�
�%�-��o���&¹��\��X�����u���d�o�;�G���������Z�����u�0�0�<�w�<�W�ԜY���F��S�D�ߊu�u�u�u���#���Y���l�N��Uʱ�;�
���w�c�D��Y���F��X��"����h�u�a�]�}�W���Ӌ��NǻN��U���<�e�h�u��%�>�������9��P1�L���u�u�u�u�3�(�W�������Z��Q��M؊�d�n�_�u�w��(�������]��1�� ���u�:�%�;�9�}�1ٚ�H����lV��G��*���&�c�
�_�w�}�����ơ�CF�N��U����u�k�d�]�}�W���Y����`2��rN��U���u�u�u�u�3�3�(���-���U��=N��U���u�:�!����J���M���F��E�����_�u�u�u�w�4�G��Y����w/��x��D���'�2�f�e�{�}�W���Yӂ��GF�
�����;�d�3�
�o��F��s���U9��Z�����d�;�
�m��h�F���Y�Ư�^��R ������b�b�
��(�(���&�Ѣ�lW��h]��D���u�2�;�'�4�0����Y���F��sN��U���u�u�u�u���$���<���JǻN��U���<�e����`�W��s���F�S��*����u�k�d�{�}�W���Yӂ��G9��s:��H���`�_�u�u�8�)����Q���F�
��E��u�
�4�g�e����Lǹ��l�N��Uʱ�;�u�k�3�'�)����K�ғ�l��h]�F�ߊu�u�u�u�8�)�J���&����lT��Q��B���%�|�_�_�]�}�W��Y����P��R �����0�}�%���.�^ϱ�Y����@��RN�����0�u�x�u�w�<�(�������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N�����
�&�u�h�6��#���H����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�&�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�e�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���#�1�%�0�w�`��������_	��T1����u�u�u�u�w�1����Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���Z ������!�9�2�6�f�`��������V��c1��Gڊ�&�
�l�|�#�8�W���Y���F�N��U���u�u�u�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���F�N�����3�}�%�&�0�?���PӒ��]FǻN��U���u�u�u�u�w�}�W���&ù��l��h����u�
�
�%�!�9�}���Y���F�N��U���0�1�<�n�w�}�W���Y���F��Y
�����u�u�u�u�w�}������ƹF�N�����3�_�u�u�9�}����
��Ɠ9F�C����%�0�u�&�>�3�������KǻN��*ڊ�'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}����	����[��G1�����9�f�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʥ�e�4�
�9�~�<�ϰ�����C9��Y�����6�d�h�4��4�(�������@��Q��E���;�u�4�
�8�.�(�������F��h�����|�|�!�0�w�}�W���Y���F�N��U���
�'�2�i�w��L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�d�4��1�(���Ӈ��Z��G�����u�x�u�u�'�l��������V��D�����:�u�u�'�4�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�r�r�w�5����Y���F���]���'�!�h�r�p�}����Y���F�N��U���
�
�%�#�3�-����DӇ��P	��C1�����e�_�u�u�w�}�W�����ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��U���%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��d�^Ϫ���ƹF�N��U���u�u�u�u�w�}�(ށ�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-�������� O��_�����u�u�u�u�w�}�W���Y���C9��V�����'�2�i�u���������F�N��U���u�u�u�0�3�4�L���Y���F�N��U���u�3�u�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=dךU���x�%�d�%�2�}����Ӗ��P��N����u�
�
�'�0�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӖ��l��PN�U���6�;�!�9�d��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����N��h�����:�<�
�u�w�-��������`2��C_�����|�4�1�}�'�>��������lV������!�|�u�;�w�<�(���
����T��N�����4�
�9�|�~�)����Y���F�N��U���u�u�
�
�%�:�K���&��ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�o��������V��D��ʥ�:�0�&�u�z�}�WϮ�K����E
��G��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�
��-����	����[��G1�����9�2�6�e�]�}�W���Y���V
��=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���<�u�}�%�4�3��������[��G1�����0�
��&�e�����@����[��=N��U���u�u�u�u�w�}�W���Y����R��[
�����i�u�%�6�9�)��������F�N��U���u�u�u�u�2�.����	����l��hY�U���;�_�u�u�w�}�W���Y���F�N��G���
�9�
�'�0�a�W���&����_��N��U���u�u�u�u�w�}������ƹF�N��U���u�u�;�u�1�}�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ_�u�u�x�'�o����Y����T��E�����x�_�u�u����������]9��X��U���6�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��R��u�=�;�u�w�}�W���Yӏ����E��H��r�u�=�;�w�}�W���Y���F��h\�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�}��������]��[����h�%�g�4��1�^�������9F�N��U���u�u�u�u�w��(������C9��=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�L����E
��G��U���<�;�%�:�2�.�W��Y����lS��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(ځ�	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ����F�N��U���u�u�u�<�w�u��������\��h_��U���&�2�6�0��	���&����_����ߊu�u�u�u�w�}�W���Y���F��1��*���
�'�2�i�w�-��������Z��d��U���u�u�u�u�w�}�Wϻ�
���R��^	�����`�u�=�;�]�}�W���Y���F�N��U���%�`�4�
�;�����E�Ƽ�9��h��N���u�u�u�u�w�}�W���YӃ����=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϮ�L����TF��D��U���6�&�{�x�]�}�W���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�'�2�i�w�-��������9��=N��U���u�u�u�9�2�}�W���Y���F���]���%�6�;�!�;�:���DӇ��P�V �����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�h���������YNךU���u�u�u�u�w�}�W���&ƹ��V�
N��@�ߊu�u�u�u�w�}�W����ƥ�FǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�}���Y����9��h(��*���%�&�'�2�c�d�����Ƽ�\��D@��X���u�<�
�<��/�;���&����T9��1�����
�'�6�o�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���F�N�����<��'��8��(���&����[��{1��*���
�:�%�d�a�/���K��ƹF�N��U���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	���&����S����ߊu�u�u�u�w�}�W���Y�ƥ�l
��q��9���
�
�0�
�b�}�JϿ�&����G9��1����u�u�u�u�w�}�W���Y����F�N��U���0�1�<�n�]�}�W���Y����Z ��N�����%�:�0�&�]�}�W��Y����T��E�����x�_�u�u�%�>��������XOǻN�����_�u�u�u�w�;�_�������E����U���6�>�h�r�p�}����Y���F�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�m�3�8�`�t�W������F�N��U���u�g�'�2�d�n�W��?����lS��h����u�u�u�u�w�}�W���7����l��h]�A��u� ����;�(��&����F�N��U���u�u��;�2���������l��E��F��u�h��;�2���������l��Q��D���%�n�u�u�w�}�W���Y����R��1�����'�&�g�<��8�(��I���a��R_�����0�:�
�
�f�;�(��O����9F�N��U���u�u�u�4�0�o��������9��h��*��m�i�u�4�0�o��������9��h��D���
�f�_�u�w�}�W���Y���Z��1����d�u�h�<�:�o����J˹��l�N��U���u�u�u�<�:�����A���F��Z�� ���m�%�n�u�w�}�W���Y�����R	��*���
�m�c�i�w�/����H����^��G_��Fʱ�"�!�u�f�l�}�W���Y���F������0�
�m�m�k�}����/����_��G_��Fʱ�"�!�u�f�l�}�W���Y���F���Gڊ�d�'�2�f�c�}�JϮ�H�֓�9��h_�G���n�u�u�u�w�}�W���YӖ��R
��1����b�u�h�%��1�(ց�����l��=N��U���u�u�u�u�w�?�F�������F���D���
�m�
�f�]�}�W���Y���F�E1��ۊ�0�
�m�g�k�}�(���H����P��G\�U���u�u�u�u�w�}��������l��h]�B��u�0�
�8�e����K����9F�N��U���u�u�u�0��0�Eց�����T�
N�����%�l�3�
�o��E�ԜY���F�N��Uʦ�9�!�%�`�%�:�D��Y����V
��Z�*���l�m�%�n�w�}�W���Y���F��Z��Dӊ�0�
�m�d�k�}����Hʹ��lQ��h����u�u�u�u�w�}�W���&����A��V�U��%��9�
��(�@���	������Y��D���_�u�u�u�w�}�W���Y����U��R	��M��i�u�8�
�d�;�(��&����F�N��U���u�u�!�%�f�/���K�����h_�� ���c�%�n�u�w�}�W���Y�����h]�����f�c�u�h�#�-�Dׁ�����l��=N��U���u�u�u�u�w�0�(�������
T��S�����l�3�
�c��o�}���Y���F�R ����u�u�u�u�2�9���Y����]��E����_�u�u�x�6�.��������@H�d��Uʥ�:�0�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��|�!�0�_�w�}�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��CW�����|�|�!�0�]�}�W���Y���F�e��ۊ�9�
�;�&�e�4����J����[��V ��D���9�:�0�
�����H����l�N��U���u�u�u��9�8�(���&����@9��^1����m�u�h��9�8�(���&����@9��^1��*��l�%�n�u�w�}�W���Y�����E��*���0�
�l�b�k�}����&¹��U��^����u�u�u�u�w�}�W�������V��Y�����f�m�u�h�3�1��������U�� V����u�u�u�u�w�}�W�������V��h\�*���0�
�l�f�k�}��������R��a1��*��f�%�n�u�w�}�W���Y�����D�����'�2�f�c�w�`��������U��V�����f�1�"�!�w�n�L���Y���F�N��U���4�g�a�'�0�n�B���DӖ��R
��1��*��`�%�n�u�w�}�W���Y�����h\�����f�b�u�h�#�-�E݁�����9��d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԜY�����^	�����0�&�u�x�w�}�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�F�������F�N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�e�;���P����[��N��U���u�u�u�u��3�ށ�����V��h��*��`�i�u�4�0�l��������9��h\�D���n�u�u�u�w�}�W���YӴ��T��V�����&�a�'�2�c�n�W��+����9��[1�����a�3�
�l�`�-�L���Y���F�N��U���2�g�4�9�8�8�(܁�����V�
N�����
�9�
�;�$�n����@�ӓ�]ǻN��U���u�u�u�u��8����J����lR��N�U���
���,�"�����	����Q��h��G���
�g�`�u�8�3���P���F�N��U���u�%��&�;��(���&����Z�Q�������!��;�4����KĹ��U��[�����c�1�"�!�w�i�L���Y���F�N��U���4�g�`�
�2��G��E�ƪ�C9��b"��:����9�<�9��o�(�������9��[����!�u�g�n�w�}�W���Y���F��h8��G���
�0�
�d�d�a�W���&����g��C1�����9�
�g�
��(�E��&��� F��@ ��U��n�u�u�u�w�}�W���Yӗ��G9��E��A��u�h�3�%�/��#�������G��N1�A���3�
�m�`�'�u�FϺ�����W�=N��U���u�u�u�u�w�?��������R��S�������,� ��(���� ����l0��B1�@ߊ�g�g�u�:�9�2�E���s���F�N��U���&�2�7�!�f�/���A��� ��h��9��� �
� �!�'�$�F���/����^��h�@���:�;�:�`�~�W�W���Y���F�N�����!�g�'�2�c�n�W������~3��N!��*���!�%�,�d�`�����A�ӓ�N��
�����`�|�_�u�w�}�W���Y���G��Z�����a�e�u�h�#�-�F�������Q��UךU���u�u�u�u�w�}����M˹��T9��[��Hʳ�%�-� ���)�:�������T��a1��*��`�%�}�f�3�*����J��ƹF�N��U���u�u�8�
�c�����H���F��G1�� ����!��9�>�1�(��&����lT��1��]��1�"�!�u�e�f�W���Y���F�N�����`�
�0�
�f�h�K�������f*��x��8���<�9�
�g�����Mƹ��S��S�����a�n�u�u�w�}�W���Y����^��Z�����d�f�i�u�:��Bہ�����
9��d��U���u�u�u�u�w�)���L����lR��N�U���
���,�"�����	����Q��h��G���
�g�`�u�8�3���P���F�N��U���u�!�%�d�a�/���O��� ��h��9��� �
� �!�'�$�F���/����^��h�G���:�;�:�g�~�W�W���Y���F�N����m�'�2�a�a�}�Jϸ�	����2��B�� ���%�,�d�b��;�(��L����R��X�����|�_�u�u�w�}�W���Y�ƹ�l��t��*��� �!�'�
�c�����I���F��h��6���
�!� �!�%��Cׁ�����9��d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԜY�����^	�����0�&�u�x�w�}�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�F�������F�N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�n�;���P����[��N��U���u�u�u�u�4��9���8����A��\��*ۊ�0�
�g�d�k�}����M�ӓ�lW��UךU���u�u�u�u�w�}����M�ӓ�lV��X�����a�a�u�h�;��(��&����BV��N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y����@��YN�����&�u�x�u�w�-����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�l�^Ϫ����F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�
�$��^�������F�N��U���u�u�3�
���8���H�ޓ�V��^�I���'�
� �a�a�-�L���Y���F�N��U���-��,� ��o�(���&����Z�P�����b�
�g�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dךU���x�4�&�2�w�/����W���F�G�����}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�I�����_�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���!�0�_�u�w�}�W���Y���Z*��C1�����!� �!�'��j�(���&����Z�^"�����&�
�!� �#�/�(��&����W��G]�U���u�u�u�u�w�}��������V9��E�� ���d�m�'�2�c�m�W������l%��R1����� �0�d�m�1��B���	��ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�w�}�Z���
������T��[���_�u�u�'�4�.�Wǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�r�r�w�5����Y���F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�a�t�W������F�N��U���u��9�
�8�����H�Г�V��\�I����9�
�:��2���O���� P��h����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���K�V�����'�6�&�{�z�W�W�������@F��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���^�Ƹ�VǻN��U���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�l�(���&���F��R ךU���u�u�u�u�w�}����&����V��R�����f�3�
�`�c�-�L���Y���F�N��U���4�g�a�
�2��G��E�Ƽ�e��hZ�����a�f�%�n�w�}�W���Y���F��R����
�0�
�e�e�a�W���&����9��h\�E���n�u�u�u�w�}�W���Yӕ��l��^�����e�l�i�u�2����&����T��G\�U���u�u�u�u�w�}��������l��hZ�A��u�0�
�8�b����M����l�N��U���u�u�u�!�'�e�(���&����Z�C��Mۊ� �g�m�
�e�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߊu�u�x�4�$�:�W�������K��N�����0�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��D���!�0�_�u�w�}�W���Y���N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�w�}�W���Y���F��A�����g�'�2�a�f�}�Jϱ�����D9��Q��A���%�n�u�u�w�}�W���Y����l0��1�*���
�l�m�i�w�����HŹ��lT��1��N���u�u�u�u�w�}�WϮ�/���� V��R	��E��i�u�
�4�e�n�(���K����CT��N��U���u�u�u�u�#�-�F�������V��S��*���g�d�
� �e�k�(��K�ƨ�D��\�N���u�u�u�u�w�}�Wϫ�����\��h ��*���
�e�l�i�w�3��������]	��Q��A���%�n�u�u�w�}�W���Y����]��Q��*؊�0�
�e�f�k�}��������9��h\�C���n�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�3�_�u�w�3�W�������9l�N�U���<�;�%�:�2�.�W��Y����A	��D�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���O��_��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���J����lW��G�����u�u�u�u�w�}�W���	����9��h��*��e�i�u�
�6�o�Bف�����9��d��U���u�u�u�u�w�-�!���&����l��hZ�A��u�
�4�g�$�o�(���J����CU��N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y����@��YN�����&�u�x�u�w�-����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�l�^Ϫ����F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�c�1�0�F���PӒ��]l�N��U���u�u�u�'�!�����K���F��AV�� ��l�
�g�_�w�}�W���Y���F�N��*����&�
�!�"�)����M˹��@��R	��G��g�1�"�!�w�t�K���;����p��h=�� ���'�
�a�
�6�)����L�ғ�N��S�����|�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǻN��Xʴ�&�2�u�'�4�.�Y��s���C��R��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������A�C�����u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���HĹ��^9��N�����-�!�:�1�1��A���	���R��X ��*���
�|�|�!�2�W�W���Y���F�N��Uʡ�%�d�a�'�0�i�E���Y����G	�N�U���
�e�
� �d�l�(��Hӂ��]��G�U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K��D��ʥ�:�0�&�u�z�}�WϮ�����N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W��PӒ��]l�N��U���u�<�u�}�6�����&����P9��
N��*���
�&�$���)�(���&����]�V�����
�:�<�
�w�}����PӇ���������7�1�d�l�~�}����Y���F�N��U���8�
�`�
�2��@��E�Ƽ�9��h��]��1�"�!�u�f�f�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߊu�u��6��<��������A��V�����'�2�a�e��}�������[�^�E��u�u�!�%�f�i����M����U��X����u�h�w�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�n�_�u�w�p��������@��RN�����
�&�|�:�w�5�W����ơ�P��R@��X���u�4�
��1�0��������\������u�4�
��1�0�W�������C9��P1����l�u�-�!�8�9����O�ԓ�OǻN�����_�u�u�u�w�<�Ͽ�&����@��Dd��U���u�u�u�"�2�}����&����U��N��U���u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Y����R��^	�����e�|�|�!�2�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����U��UךU���u�u�u�u�w�}����Y���F�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}�W�������U]ǻN��U���u�u�=�;�6��#���K����lW�	NךU���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y����[��V��!���f�3�8�g�j�}�W���Y���F�N�����
�&�u�h�6��#���M����lU��N��U���u�u�"�0�w�-�$���ǹ��^9��
P��U���u�u�u�u�w�}����*����Z�V��!���`�3�8�a�]�}�W���Y���D����&���!�
�&�
�w�c�}���Y���F�N������3�8�i�w�-�$���Ź��^9��=N��U���u�u�u�=�9�<�(���
�Г�@��S����u�u�u�u�w�}�W���7����^F���&���!�
�&�
�l�}�W���Y�����YN��*���&�b�3�8�a�`�W���Y���F�N��U����
�&�u�j�<�(���
�ޓ�@��d��U���u�u�u�"�2�}����&����U�� N��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�l�3�8�o�W�W���Y���F��R �����
�!�
�&��}�I�ԜY���F�N��Uʴ�
��3�8�k�}����&����l ��hW�U���u�u�u�u� �8�W���*����V��D��U��_�u�u�u�w�}�W���Y����`9��ZN�U����
�!�d�1�0�F��Y���F�N�����4�
��&�f�����I���9F�N��U���u�u�u�%������DӇ��`2��C_�����d�n�u�u�w�}�W�������R��c1��D؊�&�
�d�h�w�}�W���Y���F���;���&�u�h�4��	���&����T��N��U���u�u�"�0�w�-�$����Փ�@��N��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�d�
�&��n�}���Y���F�@��U����
�!�a�1�0�F���G���F�N��U���u�4�
��1�0�K���	����@��h��*��_�u�u�u�w�}�W���Ӈ��`2��C_�����d�u�k�_�w�}�W���Y���F��h �����i�u�%���)�A�������9F�N��U���u�=�;�4��	���&����S�	NךU���u�u�u�u�w�}����&����[��G1��*���b�3�8�d�l�}�W���Y�����YN��*���&�d�
�&��k�J���Y���F�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�;�!�}�/�)��������T��N�����:�&�
�#��t�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��L���8�d�n�u�w�}�W���Y�����Rd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�d�
�&��j�}���Y���F�N�����<�n�u�u�w�}�W�������R��c1��DҊ�&�
�b�h�w�}�W���Y���F���;���&�u�h�4��	���&����P��N��U���u�u�"�0�w�-�$����ߓ�@��N��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�g�
�&��d�}���Y���F�@��U����
�!�e�1�0�F���G���F�N��U���u�4�
��1�0�K���	����@��Q��E�ߊu�u�u�u�w�}��������@F�NךU���u�u�u�u�w�}����&����[�o6��-���������U�ԜY���F��SN����u�u�0�1�'�2����s���uT��h��C���%�u�h�&�3�1��������AN��D�����%�6�;�!�;�l�(��P����]��Y�����f�
� �c�g�-�^��Y����9��h[�*��i�u�!�
�8�4�(�������]��Y�����:�&�
�#�e�i�D���Y����T����*܊� �`�g�%�~�f�W���(����z(��1��*��
�g�i�u�f�}����Q����V��1�����`�
�g�u�w�4��������]��[�*��|�0�&�u�g�f�W���(����z(��Q��AҊ�g�i�u�d�w�5�������� ��Q��A؊�g�u�u�<�9�9��������_��h_�\ʰ�&�u�e�n�w�}�%���¹��_9��R��*���d�b�
�g�k�}����&����Q��G\�����8�
�g�3��h�@���P���F��Y	��*���
�;�&�g�1��G���	���N��Y	��*���
�;�&�d�>����L˹����<�����4�9�:�0�����Iǹ��]ǻN�����d�4�9�:�2��(���HĹ��lW��1��U��}�4�'�
��l����A�ԓ�F��SN�����
�9�
�;�$�o�ށ����� U�=N��U���2�d�4�9�8�8�(݁�H����W��h�I���u�u�u�u��3�ށ�����V��h��D��
�g�"�0�w�2�(�������ZW��B1�C܊�g�e�u�u�f�t����Y���F���*���f�
� �d�d��D�ԜY�ƞ�]��h��*���&�g�<�d��(�E��&���F��V��*ۊ�
�0�
�l�`�<�ό�����R
��X ��*؊�
�0�
�l�`�f�W���+����9��[1�����
�
� �d�f��D��Y���F�<�����4�9�:�0��(�F��&����[�������d�b�<�3��k�N���Q���A��N�����u�u�u�u�$�1����A����Q��h����u�4�2�d�6�1����&����K9��h��D��
�g�i�u��3�ށ�����V��h�����f�f�u�;�w�<����&����ZW��B1�Lي�g�n�u�u��3�ށ�����V��h��*��� �d�c�
�e�a�Wǌ�����R
��X ��*؊�
� �d�d��n��������lW��X��*���d�a�
�g�l�}�Wό�����R
��X ��*ي� �d�e�
�e�a�WǪ�	˹��l_��h����!�%�`�
�"�d�C���P���F��Y	��*���
�;�&�`�1��N���	���D�������
�0� �!�f�;�(��H����F��h�����#�
�|�0�$�}�G��Y����R��1�����0�
�
� �d�n�(��E���F��R �����&�9�
�
�2��F��DӇ��P	��C1��F��u�9�0�w�u�W�W�������l��h�����
�c�`�%�w�`�_����ԓ�_
��Y��D���3�
�c�d�'�}��������l��h�����3�
�`�b�'�t�}���Y����VW��[�����
�
� �d�`��E��Y���D��F�����3�
�d�`�'�}�W�������l
��1�U���0�w�w�_�w�}����H����l��X��*���d�m�
�g�k�}�%���¹��_9��R��*���d�e�
�g�/�/��������_��G�U����;�0�
�;�����&����l ��_�*��i�u�u�u�w�}���K����U��W�����=�;�}�'�4�3�F���¹��lW��1��]���h�r�r�u�;�8�}���Y���@��C��L���
�d�m�%�l�}�Wό�����R
��M�����<�3�
�b�n�-�W��s���F�G1�G���3�
�c�f�'�}����Q����\��Y��*���d�f�
�g�g�}�W��PӃ��VFǻN��U���0�
�8�d��(�F��&����F�e��ۊ�9�
�0�:�����I����Z�_�����u�8�;��a�;�(��&�����T�����`�
�|�0�$�}�G��Y����R��1�����'�&�a�3��d�@���Y���D��_��]���0� �!�d�1��N���	���R��X ��*���
�|�0�&�w�m�L���YӴ��T��V�����&�`�3�
�e�d����D������YN��*��� �!�a�'�0�i�@���Y����\��h��*���0�&�u�e�l�}�Wό�����R
��M�����
�c�b�%�w�`�_����ד�_
��Y��D���
�`�b�%�w�2�W�������l
��h_����u�4�2�g��l����O�Փ�F���*���<�
�0�!�%�.����������^	��¸�;��3�
�f�h��������G��EF�����0�}�e�u�w�0�(�������_��F�X���:�;�:�e�~�t�L���YӴ��T��a1�����e�e�%�u�j�.��������V��EF�����'�2�!� �$�:��������9��hX�*��y�:�<�!�0�/��������V�N����
� �d�f��l�D��Y����G	�G��\�ߊu�u�4�2�e�<��������U��[�����h�w�w�"�2�}�%������� 9��h_�E���u�u�
�
��(�F��&���V
��L�N���u��;�0��1�(���
�ד�9��h_�M���u�h�_�u�w�}�W����ԓ�_
��Y��D���
�e�g�%�w�5��������WW��h�����e�e�%�}�~�`�P���Y����l�N��Uʧ�#�
� �d�f��E�ԜY�ƞ�]��h��*���&�d�<�3��k�F���Y���F�N��'���0�
�9�
�9�.����O�ӓ�F��R �����:�1�d�
��(�F��&���F�_��U���0�_�u�u�w�}��������
W��UךU���4�2�g�4�;�2����&����ZW��B1�Lӊ�g�i�u��9�8�(���&����lW��1����g�u�:�u�'�>�����ד�]ǻN�����g�4�9�:�2��(���&����lW��1��U��}�4�2�g�6�1����&¹��U��]�����:�u�%�6�9�)����H��ƹF��V ��G���9�:�0�
��(�E��&���F�N�����%��&�9���N���&����l��
N��*���&�
�#�
�~�8����I��ƹF��V ��G���9�:�0�
��(�D��&���F�N�����%��&�9������H�����T�����g�f�u�9�2��U�ԜY�ƞ�]��h��*���&�3�
�c�b�-�W��[����[��<������d�3�
�a�n����Y����U��_�����0�&�u�e�l�W�W���TӇ��W	�������%�:�0�&�w�p�W�������]��D�����:�u�u�'�4�.�_�������C9��P1������&�g�
�$��N�ԜY�Ʈ�T��N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�g�;���P����[��=N��U���u�u�u�%�3�3�W������]��[����_�u�u�u�w�1��ԜY���F�N��*���0�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�1�0�6�.��������@H�d��Uʴ�
�1�0�4�$�:�(�������A	��D�����4�!�u�%�$�:����&����GW��D��\���u�7�2�;�w�}�W������]	�������!�9�2�6�f�`��������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�e�|�w�5��ԜY���F�N��*���0�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������_�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����E��ʴ�&�2�u�'�4�.�Y��s���R��R��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�o�(���&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������
O����ߊu�u�u�u�w�}�������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�'�4�.�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������
F��D��U���6�&�{�x�]�}�W���
����W��W�����;�%�:�u�w�/����Q����G��N��E���
�9�
�;�$�:�W���&����_��Y1�����
�
�%�#�3�4�(���UӖ��l��A�����<�|�u�u�5�:����Y���F�N��U���&�2�7�1�f�d�K���Q����R��[
�����2�h�4�
�8�.�(�������	����*���#�1�<�
�>�}�W�������l
��^��\ʺ�u�%�d�4��1�(���
�����T�����2�6�e�u�%�u�(߁�	����l��D��Hʴ�
�:�&�
�8�4�(�������C9��V��Hʴ�
�:�&�
�8�4�(���B����������n�_�u�u�z�}��������lW�������%�:�0�&�w�p�W�������T9��S1�L���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�d�l�i�w�<�(���
����9��
N��*���3�8�c�1� �)�W���B����������n�_�u�u�z�}��������lW�������%�:�0�&�w�p�W�������T9��S1�D���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�d�d�i�w�<�(���
����9��
N��*���3�8�b�1� �)�W���B����������n�_�u�u�z�}��������lW�������%�:�0�&�w�p�W�������T9��S1�F���&�2�
�'�4�g��������C9��h��\���u�7�2�;�w�}�W���Y���F��G1�����1�d�f�i�w�<�(���
����9��
N��*���3�8�m�1� �)�W���B����������n�_�u�u�z�}��������lT��N�����u�'�6�&�y�p�}���Y����Z��S
��D���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�g�d�w�`�_�������l
��h_��U����
�&�}�w�2����H����F�R �����0�&�_�_�w�}�ZϿ�&����Q��_�U���<�;�%�:�2�.�W��Y����C9��P1����g�
�&�<�9�-����Y����V��V��&���8�_�u�u�2�4�}���Y���F�N�����<�
�1�
�f�i�K�������]��[��D��4�
��3�:�o��������]ǻN�����'�6�&�n�]�}�W��Y����Z��S
��D��4�&�2�u�%�>���T���F��h��*���
�d�g�4�$�:�(�������A	��D�����
�&�|�u�w�?����Y���F�N��U���%�&�2�7�3�o�D���D�έ�l��D��ۊ�u�u�%���.�_�������U�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1����f�u�&�<�9�-����
���9F������7�1�g�f��.����	����	F��X��´�
��3�8�]�}�W������F�N��U���u�4�
�<��9�(��@�����T�����d�d�h�4������Mӂ��]��G����u�;�u�'�4�.�L�ԶY���F��h��*���
�d�b�4�$�:�W�������K��N�����<�
�1�
�f�j��������\������}�%��
�$�t�W�������9F�N��U���u�u�u�%�$�:����K����[�V�����
�#�
�u�w�-�4���
����W	��C��\��u�u�0�1�'�2����s���F������7�1�g�b�6�.��������@H�d��Uʴ�
�<�
�1��l�(�������A	��N�����&�4�
��1�0�}���Y����]l�N��U���u�u�u�4��4�(���&����[�V�����
�#�
�u�w�-�4���
����W	��C��\��u�u�0�1�'�2����s���F������7�1�g�b�6�.��������@H�d��Uʴ�
�<�
�1��n�(�������A	��N�����&�4�
��1�0�}���Y����]l�N��U���u�u�u�4��4�(���&����[�V�����
�#�
�u�w�-�4���
������Y��D���n�u�u�0�3�-����
��ƓF�C�����2�7�1�g�`�<����Y����V��C�U���4�
�<�
�3��B؁�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F��*���&�
�#�
�w�}����&����W��X����|�n�u�u�2�9��������9l�N�U���&�2�7�1�d�h�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&���� V��S�����:�&�
�#��}�W���:����^N��
�����d�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�n�@Ͽ�
����C��R��U���u�u�4�
�>�����HĹ��@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9�� N�U´�
�:�&�
�!��W���	����U��]�����:�d�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�D������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��\�I���4�
�:�&��+�(���Y����`9��ZF�U���;�:�d�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���HӇ��Z��G�����u�x�u�u�6���������9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�D��u�4�
�:�$��ށ�Y�ƭ�l%��Q��D���:�;�:�d�~�f�W�������A	��D����u�x�u�%�$�:����J�ƭ�@�������{�x�_�u�w�-��������9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�U��}�%��
�$�u�W������F�V�����
�#�
�|�]�}�W���Y����V��=dךU���x�4�
�<��9�(��Y����T��E�����x�_�u�u�'�.��������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h]�U��}�%�6�;�#�1�F��DӇ��p5��D��Mʱ�"�!�u�m�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����K�ƭ�@�������{�x�_�u�w�-��������T��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��G���h�}�%�6�9�)����H����C9��h��]��1�"�!�u�`�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lR��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����a�1�"�!�w�i�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��Y�����;�%�:�u�w�/����Q����`9��ZGךU���0�<�_�u�w�}�W���Y���R��^	�����a�u�h�}�'�>�����ד�[��G1��*���}�l�1�"�#�}�N���s���V��G�����_�_�u�u�z�<�(���&����R��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��Z�����;�%�:�u�w�/����Q����G��N��*���
�&�$���)�(���&����lV��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�a�i�w�u��������\��h_��U���
�%�#�1�w�3�W���Q�έ�l��D�����
�u�u�%�$�:����&����GW��D��\ʴ�1�}�%�6�9�)���������D�����|�_�u�u�9�}����
��Ɠ9F�C����<�
�1�
�d�<����Y����V��C�U���4�
�<�
�3��D���
����C��T�����&�}�%�&�6�)�W���
����@��d:��ۊ�&�
�y�%�f�<�(���P�����^ ךU���u�u�u�u�w�}��������lP��S�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�$�<����Y������T�����2�6�d�h�'�l�������9F���U���6�&�n�_�w�}�Z���	����l��hY����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1�����9�|�u�u�5�:����Y���F�N��U���&�2�7�1�`�}�J������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��G���
�9�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�O���
������T��[���_�u�u�%�$�:����Aƹ��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(ځ�	����l�N�����u�u�u�u�w�}�W�������T9��S1�U��}�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����_�d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�d�
�$��W�������A	��D�X�ߊu�u�%�&�0�>����-����9��Z1�����2�
�'�6�m�-����
ۇ��@��U
��G��_�u�u�0�>�W�W���Y�ƥ�N��h��*���
�d�|�!�2�}�W���Y���F��G1�����0�
��&�f�����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�<�
�&�&��(���I����l_�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����D�����
��&�d��.�(������]F��X�����x�u�u�4��4�(�������@��h��*���4�&�2�
�%�>�MϮ�������D�����g�b�_�u�w�8��ԜY���F��F��*���
�1�
�f�~�)����Y���F�N�����2�6�0�
��.�Fށ�
����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����9��Z1�U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C�����2�6�0�
��.�F݁�
������^	�����0�&�u�x�w�}��������V��c1��D؊�&�
�d�4�$�:�(�������A	��D�����2�7�1�g�`�W�W�������F�N�����4�
�<�
�3��B�������9F�N��U���u�%�&�2�4�8�(���
����U��_��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��C_�����d�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
����U��\�����;�%�:�0�$�}�Z���YӇ��@��T��*���&�d�
�&��o��������\������}�%�&�2�5�9�D��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���f�3�8�d�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�.��������l��1����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�f�����J����Z��G��U���'�6�&�}�'�.��������l�N�����u�u�u�u�>�}��������W9�� G�����_�u�u�u�w�}�W���
����@��d:�����3�8�d�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�a�1�0�F���DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���
����@��d:�����3�8�d�u�$�4�Ϯ�����F�=N��U���&�2�6�0��	���&����R��D�����:�u�u�'�4�.�_���
����W��Z��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��A��u�=�;�_�w�}�W���Y�ƭ�l��h�����
�!�`�3�:�l�W������]��[����_�u�u�u�w�1��ԜY���F�N��*���
�&�$���)�B�������[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�ƭ�l��h�����
�!�c�3�:�l�W�������A	��D�X�ߊu�u�%�&�0�>����-����9��Z1�*���<�;�%�:�w�}����
�έ�l��h��*��|�u�u�7�0�3�W���Y����UF��G1�����1�f�l�u�?�3�}���Y���F�V�����&�$��
�#�k����H�����T�����2�6�d�_�w�}�W������F�N��U���4�
�<�
�$�,�$����Г�@��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�V�����&�$��
�#�j����H�ƭ�@�������{�x�_�u�w�-��������`2��C_�����d�
�&�<�9�-����Y����V��V�����1�
�a�|�w�}�������F���]���&�2�7�1�d�l�W������F�N��Uʴ�
�<�
�&�&��(���N����lW��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��h��*��i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�&�&��(���A����lW��V�����'�6�&�{�z�W�W���	����l��F1��*���m�3�8�d��.����	����	F��X��´�
�<�
�1��o�^���Yӄ��ZǻN��U���3�}�%�&�0�?���K�Ƹ�V�N��U���u�u�4�
�>�����*����^��D��B��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}��������V��c1��DҊ�&�
�b�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�4�
�>�����*����_��D��Mʴ�&�2�u�'�4�.�Y��s���R��^	������
�!�l�1�0�Fׁ�
����l��TN����0�&�4�
�>�����O��ƹF��R	�����u�u�u�3��-��������S�C��U���u�u�u�u�w�<�(���&����l5��D�*���
�m�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӇ��@��T��*���&�d�
�&��e�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<�(���&����l5��D�����e�4�&�2�w�/����W���F�V�����&�$��
�#�����&����T��E��Oʥ�:�0�&�4��4�(���&���F�U�����u�u�u�<�w�<�(���&���� P�C��U���u�u�u�u�w�<�(���&����l5��D�����e�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������T9��R��!���d�3�8�e�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��h��*��4�&�2�u�%�>���T���F��h��*���$��
�!�g�;���&����T��E��Oʥ�:�0�&�4��4�(���&����9F����ߊu�u�u�u�1�u��������lR��N�����u�u�u�u�w�}��������V��c1��Gڊ�&�
�l�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�g�
�$��N��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��G���8�d�4�&�0�}����
���l�N��*���
�&�$���)�(���&¹��@��h����%�:�0�&�6���������P�N�����;�u�u�u�w�4�Wǿ�&����Q��_�\ʡ�0�u�u�u�w�}�W�������T9��R��!���g�3�8�d�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�g�1�0�F��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��F���8�g�4�&�0�}����
���l�N��*���
�&�$���)�(���&����@��h����%�:�0�&�6���������R�N�����;�u�u�u�w�4�Wǿ�&����Q��_�\ʡ�0�u�u�u�w�}�W�������T9��R��!���f�3�8�g�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�f�1�0�E��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��A���8�f�4�&�0�}����
���l�N��*���
�&�$���)�(���&����@��h����%�:�0�&�6��������� T�N�����;�u�u�u�w�4�Wǿ�&����Q��_�\ʡ�0�u�u�u�w�}�W�������T9��R��!���a�3�8�f�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�a�1�0�D��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��@���8�a�4�&�0�}����
���l�N��*���
�&�$���)�(���&ǹ��@��h����%�:�0�&�6��������� _�N�����;�u�u�u�w�4�Wǿ�&����Q��_�\ʡ�0�u�u�u�w�}�W�������T9��R��!���`�3�8�a�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�`�1�0�C��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��C���8�`�4�&�0�}����
���l�N��*���
�&�$���)�(���&ƹ��@��h����%�:�0�&�6���������Q�N�����;�u�u�u�w�4�Wǿ�&����Q��_�\ʡ�0�u�u�u�w�}�W�������T9��R��!���c�3�8�`�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�c�1�0�B��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��B���8�c�4�&�0�}����
���l�N��*���
�&�$���)�(���&Ź��@��h����%�:�0�&�6���������
OǻN�����_�u�u�u�w�;�_���
����W��W�����u�u�u�u�w�}�WϿ�&����P��h=�����3�8�c�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�b�3�:�k�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�<�(���&����l5��D�����b�4�&�2�w�/����W���F�V�����&�$��
�#�����&����T��E��Oʥ�:�0�&�4��4�(���&����9F����ߊu�u�u�u�1�u��������lW��N�����u�u�u�u�w�}��������V��c1��M���8�b�i�u�'�>��������lW��N��U���0�&�u�u�w�}�W���YӇ��@��T��*���&�m�3�8�`�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����
����g9��1����4�&�2�u�%�>���T���F��h��*���$��
�!��.�(ׁ�
����l��TN����0�&�4�
�>�����@��ƹF��R	�����u�u�u�3��-��������
U�C��U���u�u�u�u�w�<�(���&����l5��D�����m�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������T9��R��!���l�3�8�m�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R�����u�7�:�
��m��������A9��h+�����
� �g�e��o�K�������U��B1�Eڊ�f�-�'�4��2����¹��l�N������e� �
�%�<��������R
��h��G���
�g�i�u�#�-�F�������V��O�����:�&�
�#��t�}���Y����l��N!��*���4�0�
�'��(��������V��N�U �!�3�
�`�c�-�W���Y����\��h��*���_�u�u�'�2�:�F�������T��^_�� ��l�
�g�i�w�3� �������9��h_�M���u�;�u�0�2�8�(���
�֓�9��h_�M���|�_�u�u�%�8���H����\��Y1�����d�`�%�u�j�u��������l��h]�Fʴ�1�1�9�!�3�2����&����lT��1��\�ߊu�u�'�0�0�l�F���&����V��G\��H���'�0�2�d�f�9��������l ��W�*��-�'�4�
�8�.�(���&����F�U�����g�
�
� �e�e�(��E����A��P�D���8�'�4�
��(�E��&����\��G1�����9�d�d�n�w�}�������� 9��h��D��
�g�i�u�4�/��������9��h_�F���u�'��;�2���������l��h�����m�l�%�|�]�}�W�������U��h��D��
�g�i�u�4�/��������l ��Y�*��:�u�4�2�e�<��������]	��^1��*��`�%�|�_�w�}�����ד�F9��_��G��u�!�%�d�1��G���	�ƣ���R��D���1�8�'�4��l����@�ӓ�O��N�����'�0�e�1�:�/����H���� W��h�I���;�"�<�;�>��(���J����CU��Y
�����0�
�;�&�e�;�(��O����l�N�����0�e�1�8�%�<�(�������V��N�U»�"�<�;�<�����Hù����
�����
�;�&�f�1��E���	����F�U�����e�1�8�'�6��(���K����CT�
N�����<�
� �g�o��DϿ�ӈ��@��U��G���
�f�c�%�~�W�W�������V9��h\�E���u�h�}�8�b�;�(��M����\��E����d�1�8�'�6��(���K����CT�=N��U���0�2�
�d�1��N���	���N��@�����
�
� �d�a��Dϱ�Y����G��M�����;�!�<�
�"�l�@܁�K��ƹF��E�����g�3�
�a�e�-�W��Q����Z��^��*���g�`�
�f�8�}�(���&����lT��1��\�ߊu�u�'�0�0��D���&����l��S�����<�;�<�
��(�D��&����AF��Y��ۊ� �f�l�
�e�f�W�������T��1��*��f�%�u�h��8��������l ��\�*��:�u�
�:��o����K�ѓ�O��N�����'�0�<�3��l�N���Y���]��^	�����0�
�l�f�8�}��������A	��1�����3�
�d�a�'�t�}���Y����A��^1��*���g�d�
�g�k�}��������lW��B1�E݊�g�:�u�#�%�1� �������_��G�U���7�8�'�0�>�4�(���K����CT�
N�����3�:�
�
�2��G���ƣ�V��X��*���
�e�m�n�w�}��������l��Q��D���%�u�h�}�9�8����&����lU��1��U���:�0�3�:�����Hƹ��]ǻN�����2�
�
�a�1��D���	���N��S�����a�3�
�f�o�-�W�������_	��1��*��a�%�|�_�w�}��������Z9��h\�G���u�h�}�;�2�;��������9�������3�:�
� �e�k�(��B�����h^��G���4�1�0�&�w�`����H�ғ�F9��Z��D��x�d�1�"�#�}�^�ԶY���F��Q1��D��
�1�'�&�f�<����Y����V��C�U���7�3�e�d�c�����
�ד�@��Y1�����u�'�6�&��-��������`2��C_�����d�y�4�
�>�����*����P��D��@���%�&�2�6�2��#���Hƹ��^9��d��Uʷ�2�;�u�u�w�}����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y����9��W�����&�d�i�u�'�>��������N��N����!�u�|�_�w�}�W�������N��h�����:�<�
�u�w�-��������`2��C_�����d�|�u�=�9�W�W���Y���F��Q1��D��
�1�'�&�f�a�W�������l
��1�G���d�1�"�!�w�t�}���Y���V
��QN�����:�&�
�:�>��W���	����l��F1��*���a�3�8�d�~�}����s���F�N�����e�d�a�
�3�/���E�ƭ�l��D�����e�g�x�d�3�*����P���F�N�����u�u�u�u�w�}����I����
9��S�����h�w��n�w�}�W�������U]�N�����%�:�0�&�]�W�W���Tӄ��lV��Z����4�&�2�u�%�>���T���F��Q1��D��
�0�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
����U��X��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����Q��D��C���u�=�;�_�w�}�W���Y�Ʈ�U9��\�*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W�������T��h��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C�� ���
�g�l�6�f�<����Y����V��C�U���7�3�e�d�c��ށ�
����l��TN����0�&�4�
�2�}��������B9��h��A���8�d�y�4��4�(�������@��h��*���u�%�&�2�4�8�(���
����U��Z��U���7�2�;�u�w�}�WϷ�Y���R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���u�'�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�a�;���P�ƣ�N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��[�����a�|�|�!�2�}�W���Y���F��B��*��l�6�d�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����F ��h_�L���d�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���7�3�e�d�c��FϿ�
����C��R��U���u�u�7�3�g�l�Cց�H����Z��G��U���'�6�&�}��>�(�������F��E��Bۊ�0�
�d�c�w�-��������`2��C_�����d�y�<�
�#���������F��Y�����a�e�y�4��4�(�������@��h��*���u�%�&�2�4�8�(���
����U��Z����!��&�
�#�(����&����U��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w�-��������`2��C_�����d�|�u�=�9�W�W���Y���F��Q1��D��
�d�i�u��>�(�������F��E��Bۊ�0�
�d�c�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��@���8�d�|�u�?�3�}���Y���F�U��E��a�
�d�i�w���������G��C��*��
�0�
�g�f�W�W���Y�Ʃ�@��F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�5��ԜY���F�N�����d�a�
�d�k�}�;���&����l5��B�����m�
� �f�o��D�ԜY���F��D��U���u�u�u�u�5�;�G��Mʹ��Z�6��-���������/���!����k>��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u� ���E�������@��YN�����&�u�x�u�w�?����H����D��V�����'�6�o�%�8�8�ǿ�&���R��^	������
�!�a�1�0�F������T9��R��!���d�
�&�
�b�}��������B9��h��@���8�d�|�u�w�?����Y���F��QN��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���a�3�8�d�~�}��������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����Г�@��G�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��i�^�������9F�N��U���u� �
�
�e�d� ��E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���
�
�g�l� �l�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�u�u�6�%�$�F���&����l��S�����d�m�'�2�c�m�W���Y����
W��B1�@ӊ�g�n�u�u�4�/����¹��lW��1��U��}�0�
�8�d����HŹ������B���
�m�c�%�~�W�W�������9��Q��@���%�u�h�}�2���������V��N��ʡ�%�
� �d�n��E��Y����R��h_�����d�3�
�m�d�-�W��Q����l ��V�*��:�u�8�
�e����I˹��]ǻN�����
�
�:�
��(�F��&���F��Z�����b�f�%�u�%�)���&����W��G]����u�4�'�
��(�D��&���F��Z��@ߊ�0�
�d�m�6�9����@ƹ��lU��1��\�ߊu�u�4�'��(�E��&���F��Z��Aڊ� �g�g�
�d�<�Ϫ�	����U��X�����_�u�u�0�2�8�(���
�֓�9��h_�M���u�h�}�0�2�8�(���
�ד�F9��[��Fʺ�u�0�
�8�c����J����]ǻN�����0�
�;�&�g�4����H�ד�F�F�����1�:�0�
�2��N���ƿ�_9��G\�����d�c�%�|�]�}�W�������\��h_�� ��d�
�f�i�w�}�W���YӴ��T��V�����
�
� �
�f�;�(��I����D��F�����0�g�
�d�1��N���	����[�I�����u�u�u�u�w�-�F���¹��T9��[�U���1�9�!�1�8�8�(݁�����9��R�����u�u�u�
�f�4�(���J����CT��_��]���'�
�
� �d�k�(��I���W����ߊu�u�u�u�6�:�F�������@9��E��A��n�u�u�1�;�)��������U��X�����h�_�u�u�w�}�(�������lU�� 1��U���;�}�4�'�����Kǹ��V�
N��R���9�0�_�u�w�}�W����ד�_
��Y��C���
�g�a�%�l�}�WϺ�����l	��D1��*��b�%�u�h�]�}�W���Y����VW��[�����g�8�-�<�1��@���	�ƻ�V�U�����g�
�
� �f�k�(��I���W����ߊu�u�u�u��o�(�������9��d��Uʱ�9�!�1�/�%�.�G�������U��Y�����h�}�8�
�n�/���K�ƭ�WF��[�����'�&�d�;�#�;�(��N����l�N�����1�/�'�&�g�3��������R��N�U¡�%�g�
�0��d�GϿ�ӂ��V��h�����:�
� �g�c��E��Y����V
��R
�����
�
� �d�`��D��Y���F�<�����4�9�:�0���F������� F��R �����,�d�<�
�"�l�A݁�K���F�G�����_�u�u�u�w�<��������V��h\��D���2�f�a�n�w�}��������V��h_����� �d�c�
�e�a�WǺ�����l��X��*���d�b�
�f�/�/��������_��G�U���1�9�!�1�-�/��������^��N�U¦�2�7�!�3��o�O���Y����]	��T�����
�f�g�%�~�W�W�������W9��E��F���
�e�e�%�w�`�}���Y���a��R_�����;�&�`�'�0�i�E������P��N1�����e�`�%�}�~�`�P���Y����l�N��Uʇ�;�0�
�9��8����&����W��d��Uʱ�9�!�1�/�%�.�C���&����l��S��U���u�u��;�2���������l ��\�*��"�0�u�6�%�$�E���&����l��G��U��|�0�&�u�w�}�W���+����9��[1�����`�3�
�g�n�-�L���Yӂ��V��h����� �g�e�
�d�a�W���Y���4��P�����:�0�
�
��8�(��Nӑ��]F��V��*ۊ�
�0�
�l�`�m�W���H����_��=N��U���u�4�2�d�6�1����
�ԓ�l��h]�F�ߊu�u�0�0�2�����&����U��Z�����h�}�0�0�2�����&����V��G]�����%�6�;�!�;�l�F��Y����K��X �����c�g�%�u�j��Uϩ�����9��h(��*���%�&�'�2�c�d�JϿ�&����G9��1�U���0�w�w�_�w�}����&¹��lP��h�I���!�
�:�<��8����
����WN��h�����#�g��d�w�}����ے��lU��Q��Dڊ�d�|�_�u�w�%�(�������l��S�����:�<�
�0�#�/�����έ�l��D������d�u�u�>�3�Ǫ�	�Г�F9��1��\��u�u�0�%�#�-�!�������9��R�����
�
�
� �b�i����Kӂ��]��\����u�-�
�8�����K����[��E��#���
�l�
�d�a�}��������l�N�������!��$�1��������
Q��h��G��
�f�i�u�w�}�W���	����9��h��*��m�"�0�u�#�-�@܁�����
9��^��H��r�u�9�0�]�}�W���Y����r$��x��4���9�!�
�4�"��@�������R��UךU���-�
��-�"���������R
��hW�����
�a�a�%�w�`��������l��C�� ���2�0�}�%�4�3����Kǹ��K��Y�����%��9�
�a�/���@���9F���*���-� �
�7�8�(��������
9��Q��@���%�u�h�_�w�}�W���&����lR��Q��A���%�u�=�;��0�(�������R��F�U���d�|�0�&�w�}�W���YӀ��l'��O!��*���:� �0��;�8�Nց�&����T��G\�U���3�%����)�6�������e��R1�*��� �g�g�
�e�a�W���&����P9��T��]���<�;�1�4��2�����ғ�F�B �����}�
�4�g�c����@����O��N�����;�1�
�0�:�i�@�������W��N�U���
�:�<�
�2�)�ǫ�
����WN��h�����#�`�e�u�w�3����ۀ��l��R1�����a�
�
� �e�i�(��P���F��G1�����0�8�`�d��;�(��I����[��C
�����
�0�!�'�"�.����Q����\��h��@��u�u�;�<�9�9��������G��h[�*��� �g�`�
�f�t�}���Y���U��Y��*���8�`�c��1��A���	�����h�����0�!�'�'�$�'�_�������l0��1�*���
�e�a�y�b�t�}���Y��� ��h �����'�
�a�
��(�E��&���F��S1�����#�6�:�}�2�4�ǭ�����C9��[\��C���2�f�l�|�e�t�L�ԜY�ƪ�C9��E��G����3�
�e�d�-�W��s���F�G1��؊�e�8�-�3��m�@���Y����N��[1�����3�
�e�m�'�u�^��^���V
��d��U���u�&�9�!�'�i����I�ߓ� ]ǻN�������,� ��(���� ����l0��B1�Aߊ�e�i�u�8��e����A�ԓ�N��C��U���;�:�e�n�w�}��������J)��h#�����,�d�a��1��O���	�����hZ�� ��d�
�g�_�w�}����4����|��z�����
�g�
�
�"�o�Cځ�K���@��[�����6�:�}�0�>�8��������@��[�����6�:�}�<�9�9��������J)��h#�����,�d�a��1��O���	�����Y�����-� ���#���������9��Q��M���%�|�|�u�`�t�}���Y����K+��c�����9�<�9�
�e��(���K����CV�
N����
� �g�a��l�D���Y�ƨ�D��^����u�-�
���$��������_��Y��*���g�`�
�d�k�}�(���&����U��G\�U���3�%�-� ����������J9�� 1�����m�`�%�u�j�.��������V��EF�����}�;�<�;�3�.��������V��EF�����}�-�
���$��������_��Y��*���g�`�
�e�w�}����ۀ��l��{:�� ��� �!�%�,�f�j�!���&����l��G�@���n�_�u�u�z�:����&����P��D��ʥ�:�0�&�u�z�}�WϹ�	����Q��T�����;�%�:�u�w�/����Q����Z��D��&���!�
�&�
�{�<�(���Y����Z��S
��E���4�
�<�
�$�,�$���Ĺ��^9�������6�0�
��$�o����H�ƭ�l��h�����
�!�
�&��q��������V��c1��A���8�f�u�%�$�:����&����GS��D��Yʴ�
�<�
�&�&��(���&����OǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9�_���	����@��X	��*���u�%�&�2�4�8�(���
�ד�@��N��ʻ�!�4�
�<��9�(��P�ƣ�N��h�����:�<�
�u�w�-��������`2��CY�����|�:�u�4��2��������F�V�����&�$��
�#�����PӉ����T�����2�6�d�h�6�����
����g9��1����u�'�}�%�4�3��������[��G1�����0�
��&�c�;���Y���R��X ��*���<�
�u�u�'�.��������l��h��*���:�u�4�
�8�.�(�������F��h��*���$��
�!��.�(���P�Ƹ�V�N��U���u�u�2�%�1��@߁����R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���'�
� �a�g�>�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������l��V�����'�6�&�{�z�W�W�������lR��h�����2�
�'�6�m�-����
ۇ��@��T��*���&�d�3�8�g�}����UӇ��@��U
��D��u�%�&�2�4�8�(���
�ѓ�@��N��*���
�&�$���)�(���&����C9��P1������&�f�3�:�o�W���
����@��d:��ފ�&�
�y�4��4�(�������@��Q��A���%�&�2�6�2��#���O����lS�N�����;�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�W�������]��[����h�4�
�<��.����&����U��G�����:�}�%�&�0�?���@����AF��G1�����9�2�6�d�j�<�(���&����l5��D�����c�u�'�}�'�>��������lW������6�0�
��$�o����H�ƣ�N��h�����:�<�
�u�w�-��������`2��C]�����|�:�u�4��2��������F�V�����&�$��
�#�����PӉ����T�����2�6�d�h�6�����
����g9��1����u�'�}�%�4�3��������[��G1�����0�
��&�a�;���P����[��=N��U���u�u�u�'��(�C��������T�����2�6�d�_�w�}�W������F�N��U���2�%�3�
�`����Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�>�����
����A��B��D���a�3�
�f�o�-�W��
����\��h�����&�2�0�}��>�(�������F��E��BҊ�
� �f�m��l�W���������V����
�0�
�d�c�t�}���Y����G9��D�����!�'�
�b��(�D��&���FǻN��U���0��9�d�1��B���	�ƻ�V�X�����
� �f�e��o�G���Y�����RNךU���u�u�0��;�m����M�ғ� ]ǻN��U����6�
�4�2���������^��h��F��
�d�i�u�#�����&����\��R��¦�2�0�}�8��e����J�ғ�O�G����u�<�
�!��.�(�������V9��1��*���a�%�u�h�]�}�W���Y����V
��h��F��
�f�"�0�w�2�(���ƹ��lU��1��]���h�r�r�u�;�8�}���Y���]��R�*���f�f�
�f�]�}�W�������@��C�����
�m�
�
�"�n�N܁�K���@��[�����6�:�}�;�>�3�Ƿ�&����R��d�����0�d�d�a�1��D���	�����^	��¥��9�
�c�%�:�C��P��ƹF��{1��*���0��'�6�"�8�F�������S��N�U���u�u�u�;� �8�Fׁ�����9�������'�6�;�`�1��B���	����[�I�����u�u�u�u�w�3� ���HĹ��lU��1��N���u�<�
�<��/�;���&����U��^�����h�&�1�9�0�>�����ι�@��R
��9���
�:�
�:�'�.����M���F��D�����%�6�;�!�;�o�F���s���Z*��X
�����
�f�
� �d�k�(��E�ƿ�W9��P�����:�}�;�<�9�9����A���� U��h�U���;�<�;�1�'��݁�&�ד�V��V�\�ߊu�u��!�%�l�>�������R��t�����
� �f�e��n�K���Y���F��G1�����9�f�
�u�?�3�_���&����l ��Y�*��e�u�u�d�~�8����Y���F��R�����3�
�c�f�'�f�W���Y����9��b"�����
�d�
� �d�o�(��E�ƿ�W9��P�����:�}�0�<�2�.����Q����V��Q��B���%�|�f�|�l�W�W���5����q��C1�L���
�b�f�%�w�`��������l��C�� ���2�0�}�
��3����Y�ƹ�@��R
��9���'�d��
�6�:�(���&����P��h��F��
�f�|�_�w�}����&����T��N�U��u�=�;�}�>�3�Ǫ�	����l ��W�����i�&�2�0��-��������lW������w�_�u�u�4�-�(���@�ޓ�F�L�U���;�}�<�;�3�)���I����
T��GZ��Kʦ�2�0�}�%�4�3����H¹��F��D��E��u�u�<�8�d���������9��R��]���%�
� �g�a��EϦ�Ӈ��P	��C1��D��n�u�u�<�:�n����L�ғ�F�L�U���;�}�8�
�c����LŹ��[��G1�����9�g�e�u�;�8�U���s���Z��h��@���%�u�h�w�u�*����
����WN��G1�*���`�m�%�|�i�.����Q����\��h��D��|�0�&�u�g�f�W�������e9��Q��Mފ�d�i�u�
�$�4��������9��d��Uʼ�0�
�
� �c�k����Dӂ��@��Y1��*��
�d�_�u�w�.����&����
T��N�U���2��d�3��e�(��O�ƨ�D��X�N���u�9�
�
�"�d�C���Y����^��1��*��
�g�d�x�f�9� ���Y����F�[*�� ��c�
�d�i�w�0�(�������W��F�X��1�"�!�u�~�W�W���T�Ơ�lV��[��*ڊ�1�'�&�e�6�.��������@H�d��Uʹ�
�
�a�
������
�֓�@��Y1�����u�'�6�&��-��������`2��C_�����d�y�4�
�>�����*����_��D��M�ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�6�����
����g9��W�����m�|�!�0�w�}�W���Y���
��1�@���e�4�1�0�$�}�JϿ�&����G9��Z��]���u�u�:�;�8�m�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�a�t����Y���F�N��U���e�a�`�0�g�<����
�����T�����c�
�}�u�w�}�������9F�N��U���0�_�u�u�w�}�W����֓�S��h^�����&�e�i�u���}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h^��Aߊ�
�
�1�'�$�l�����Ƽ�\��D@��X���u�9�
�
�c��(߁�����@W��D�����:�u�u�'�4�.�_���&����A��\�Yʴ�
�<�
�&�&��(���@����lW�������6�0�
��$�l�(���&���F�U�����u�u�u�<�w�u��������\��h_��U���&�2�6�0��	���&����Q����ߊu�u�u�u�w�}����M�ӓ�lV��S
����i�u�8�
�g�����K���K�
�����e�n�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��h��*��|�!�0�u�w�}�W���Y����G9��Z�����4�1�0�&�w�`��������_��h\��U���u�:�;�:�g�f�W���Y����_��=N��U���u�u�u�!�g�i�B���I����A��N�Uȍ�w�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���I����l��h��U���<�;�%�:�2�.�W��Y����G9��Z�����6�e�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����ѓ�@��B�����2�6�0�
��.�Fց�
����l�N�����u�u�u�u�>�}�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���HĹ��^9��G�����4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�l�3�8�f�t�^������F�N��U���9�
�
�a���(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʹ�
�
�a�
������DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���I����l��h��U���<�;�%�:�2�.�W��Y����G9��Z�����6�d�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����ߓ�@��B�����2�6�0�
��.�Fׁ�
����l�N�����u�u�u�u�>�}�_���	����@��X	��*���u�%�6�|�6�9�_�������l
��^��U���%�&�2�6�2��#���Hʹ��^9��G�����4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�m�3�8�f�t�^������F�N��U���9�
�
�a���(���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʹ�
�
�a�
������DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�)�G��L����l��S�����e�
� �f�f��C�ԶY���F��h^��Aߊ�
�
�0�u�$�4�Ϯ�����F�=N��U���e�a�`�0�g�*�F���
����C��T�����&�}�%�6�{�<�(���&����l5��D�*���
�b�_�u�w�8��ԜY���F��F��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�b�~�t����Y���F�N��U���e�a�`�0�g�*�F��Y����\��h�����n�u�u�u�w�8����Y���F�N�����a�`�0�e� �l�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�1�(߁�Mƹ��9��S�����&�<�;�%�8�8����T���
��1�@���d�4�1�0�$���������PF��G�����4�
�<�
�$�,�$����ѓ�@��B�����2�6�0�
��.�Fց�
����l�N�����u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���Hʹ��^9��G�����_�u�u�u�w�}�W���I����l��h�����e�i�u�%�4�3����Oǹ��F�N�����u�|�_�u�w�}�W������R��X ��*���<�
�u�u�'�.��������l�� 1����|�u�=�;�]�}�W���Y���_��hZ�*���
�1�'�&�g�a�W�������l
��1�G���d�1�"�!�w�t�}���Y���V
��d��U���u�u�u�9���Cځ�&¹��W��D^��H����n�u�u�w�}�������F�R �����0�&�_�_�w�}�Zϲ�&ù��9��1�����&�u�&�<�9�-����
���9F���E��`�0�d�4�3�8�ށ�
����l��TN����0�&�!�%�f�i����M������D�����
��&�d��.�(��Y����Z��D��&���!�m�3�8�f�t�W�������9F�N��U���}�4�
�:�$�����&���R��^	������
�!�m�1�0�F���Y����l�N��U���u�9�
�
�c��(ށ�����@W�
N����a�'�2�a�e�u�W���Y����G	�UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	���&����^����ߊu�u�u�u�w�}����M�ӓ�lW��S
����i�u�%�6�9�)���&����F��S�����|�_�u�u�w�}����s���F�N�����
�a�
�
��9����H���>��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�9�
��i�(���&����R��P �����&�{�x�_�w�}����M�ӓ�lW��R^�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�f�����O�ƭ�l��h�����
�!�l�3�:�l�^���Yӄ��ZǻN��U���3�}�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�`�;���P�ƣ�N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��W�����m�|�|�!�2�}�W���Y���F��C1��A���0�d�6�e�k�}��������\��h_�U���u�u�0�&�w�}�W���Y���
��1�@���d�6�e�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�9�
��i�(���&����R��P �����&�{�x�_�w�}����M�ӓ�lW��R_�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�f�����A�ƭ�l��h�����
�!�m�3�:�l�^���Yӄ��ZǻN��U���3�}�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�n�;���P�ƣ�N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��V�����b�|�|�!�2�}�W���Y���F��C1��A���0�d�6�d�k�}��������\��h_�U���u�u�0�&�w�}�W���Y���
��1�@���d�6�d�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���9�
�
�a���(��E�ƿ�W9��P�����:�}�<�;�3�4�(���5�Ԣ�F��\�� ��g�
�d�u�w�4��������A��~ �����
�;�
�:�%�8�E���&����l��UװU���x�u�!�e�c�h��������@��YN�����&�u�x�u�w�1�(߁�Mƹ��9��1�����
�'�6�o�'�2��������F��h��*���$��
�!�o�;���P�����^ ךU���u�u�3�}��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�O�������O�C��U���u�u�u�u�w�1�(߁�Mƹ��9��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�;��(��&����D��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԜY�ơ�]9��1��*��l�%�u�h�$�9��������G	��B �����}�%�6�;�#�1�Bہ�P����]��Y�����&�9�
�
�"�l�Oځ�H����F�Z��#���3�
�f�
�e�a�W���&����P9��T��]���<�;�1�4��2�����ғ�F�B �����}�
�0� �#�j����J����O��N������c�3�
�c��D��Y���F���*���
� �c�c�'�}����Q����T9��Q��L؊�f�e�u�u�f�t����Y���F������!�b�3�
�d��F�ԜY�ơ�]9��Q��D���%�u�h�_�w�}�W�������9��h_�L���u�=�;�}�$�8�(���&����V�
N��R���9�0�_�u�w�}�W�������lP��B1�Mߊ�d�_�u�u�2���������
R��N�U���u�u�u�<��)�4���&����P��R1�D���3�
�f�m�'�}����Q����G��1����c�}�|�h�p�z�W������F�N��*����&�
�!�"�)����Aƹ��U��W����u�u�;�"�2�l�(���J����CU�
NךU���u�u�0��;����OŹ����YN�����;�f�3�
�c�i����P���A�R��U���u�u�u�;� �8�O���&����l��=N��U����9�g�3��h�D���Y���F�N�����!��&�
�#�(����&����9��h]�F���u�=�;�}�2����&����P��G\��\��r�r�u�9�2�W�W���Y�ƥ�l��t��*��� �!�'�
�`��(���J����CT��N�����0�d�
� �d�n�(��E��ƹF�N��9���
�4�0��%�>����H�ޓ�l ��]�*��"�0�u�&�;�)��������R��F�U���d�|�0�&�w�}�W���Yӏ��P��V��&���6� �0�d�b�i����J�Փ�]ǻN�����9�a�3�
�b�d����D���F�N��*����&�
�!�"�)����N˹��U��V�����=�;�}�0��0�B݁�����R�N��R��u�9�0�_�w�}�W���5����p��h=�� ���'�
�b�
��(�D��&����F�Y����
� �f�a��n�K���Y���F��R�����3�
�`�f�'�}����Q����\��h��F��
�g�e�u�w�l�^ϻ�
��ƹF�N�����9�f�3�
�b�l���Y����V��[_�����`�g�%�u�j�W�W���Y�ƥ�l��t��*��� �!�'�
�`��(���J����CW��_��]���
�8�c�
�"�n�A߁�K���F�G�����_�u�u�u�w���������G��C��*��
�
� �f�n��E�ԜY�Ƣ�D5��Y�� ��b�
�f�i�w�}�W���Yӏ��P��V��&���6� �0�d�b�i����J�Փ�F��R �����!�%�g�'�0�i�A���P���A�R��U���u�u�u�<��)�4���&����P��R1�M���3�
�f�a�'�f�W�������_W��Q��@���%�u�h�_�w�}�W�������P��B1�C؊�f�"�0�u�8�����&����Q��G\��\��r�r�u�9�2�W�W���Y�ƥ�l��t��*��� �!�'�
�`��(���J����CT��N�����0�d�3�
�a�e����D���F�N�����1�
�0�8�b�l�!���&����l��@��Uº�
�:�1�3��k�D���Q���A��N�����u�u�u�u�9�*��������9��d��Uʻ�"�0�g�3��j�@���Y���F�N�����;�1�
�0�:�h�G�������^��N�����!�%�m�
�2��G��I���W����ߊu�u�u�u�/���������V��a1��*��e�%�n�u�w�}�Wϰ�����R��V�����b�f�%�u�j�.��������V��EF�����}�<�;�1�9�*��������^��G�@���_�u�u�;� �8�D���&����l��S��U���u�u�3�%�9�9�(�������l0��B1�@ۊ�g�"�0�u�$�1����K����lR��F�U���d�|�0�&�w�}�W���YӀ��l��R1�����e�
�
� �e�k�(��s���]��R�����b�b�%�u�j�W�W���Y�ƪ�C9��S�����`�c��3��k�@���Y����N��G1�*���
�e�`�e�w�}�F�������9F�N��U���
�:�0�!�%��N؁�&����S��G\�U���;�"�0�`�1��@���	���l�N��Uʻ�"�0�f�3��j�G���Y����N��h�����
�c�f�%��t�J���^�Ʃ�@�N��U���3�%�;�1��8���I����F9��V��D�ߊu�u�0��;����Oǹ��Z�=N��U���u�0��9�e���������U��N�����:�
�:�1�1��A���	����[�I�����u�u�u�u�w�;��������A��Y��*���g�`�
�g�]�}�W���*����U��X�����h�_�u�u�w�}�;���&����l5��B�����b�
�
� �d�e�(��������h��Cۊ� �f�c�
�e�m�W���H����_��=N��U���u��6�
�6�8�$�������lW��hZ�� ��m�
�d�_�w�}����˹��lU��1��U��_�u�u�u�w���������G��C��*��
�
� �f�n��Eϩ�����V
��Z�*���f�g�
�g�g�}�W��PӃ��VFǻN��U����6�
�4�2���������^��h��F��
�d�_�u�w�8�$���&����R��G]��H�ߊu�u�u�u��<�E��&����V�������0�
�8�`��8�(��M���F�G�����_�u�u�u�w�����HŹ��T9��V�U���;�"�0�
�"�o�@؁�J���9F�N��U���
�:�0�!�%��Gف�&����S��G_�����}�0�
�8�c�����I���F�_��U���0�_�u�u�w�}��������V��^��#���
�c�e�%�l�}�Wϰ�����Q��1��*��m�%�u�h�'��݁�@����^��h�D���:�;�:�d�~�W�W�������]��h\�� ��`�
�f�i�w�����Jù��lT��1��]��1�"�!�u�d�f�W�������T��C1�����e�d�%�u�j�-�!���&�ד�F9��X��G��u�:�;�:�d�t�}���Y����Z��^��*���f�d�
�f�k�}�(���K����U��^�����d�1�"�!�w�l�L���Yӈ��l��E�� ��m�
�g�i�w�3� �������9��h\�C���u�'�%��$�1�(�������F9�� X��G��u�u�:�
�8�9�Fځ�H����V��h�I���!�%�c�
�"�l�Eہ�KӇ����1��*��m�%�|�_�w�}��������l��B1�Eي�g�i�u�!�'�o�(���H����CT��Y
�����3�
�`�d�'�t�}���Y����\��Y��D���
�e�c�%�w�`�_���&�ғ�F9��Z��Gʴ�1�'�#�
�"�d�O���P���F��h����
�
� �d�d��E��Yے��lT��Q��@���%�u�;�u�2����L¹��]ǻN�����;�d�3�
�a�i����D�ο�_9��GZ�����a�`�u�'�>�0�D�������O��N�����:�1�
� �e�d�(��E����A9��Y
�� ��b�
�g�:�w�/����H����P��h�N���u�:�
�:�3����Nǹ��Z���*���c�
� �f�a��Eϱ�Y����G��1��*��g�%�|�_�w�}�����ғ�F9��V��G��u�&�9�!�'�j����M�ғ�F����*���3�
�f�m�'�t�}���Y����\��h��F��
�g�i�u�8�����&����Q��G\��ʺ�
�:�1�
�"�n�Oׁ�K��ƹF��E1����� �g�b�
�e�a�Wǭ�����T��R	��E��:�u�0�
�:�h�(���&����]ǻN�����9�"�d�3��d�N���Y���Q��E	��ۊ� �d�b�
�e�<�Ϫ�	����U��V�����_�u�u�#�%�1� �������^��N�U·�8�'�0�<��(�E��&����]��Z��C���
�f�a�%�~�W�W�������\��h��F��
�g�i�u�5�0��������lU��1��U���u�8�
�f�1��F���	����F�X�����
�
� �f�n��E��Yۄ��V��h�����g�f�%�u�9�}����N���� T��h�N���u�:�0�3�8����Oʹ��Z������
�
� �g�b��EϿ�Ӓ��lU��Q��D���%�|�_�u�w�p�W���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��V�����;�&�2�4�$�:�(�������A	��D��*ڊ�%�#�1�u����������TOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�e�4�
�;�t�W������F�N��Uʥ�e�4�
�9��3����E�Ƽ�9��h��N���u�u�u�0�$�}�W���Y���F��h^�����1�<�
�<�w�`��������W9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�g�4�(���Y����T��E�����x�_�u�u����������Z��G��U���'�6�&�}��q����	������h�����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�-�G���&����F��R ��U���u�u�u�u�'�m���������d��U���u�0�&�u�w�}�W���Y����lV��Y1����u�
�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����
9��h��D��
�g�i�u��3�ށ�����A	��1��*��g�%�u�'�%�+�(���@�ޓ�O��N����l�<�3�
�a�l����D�Ξ�]��h��*���:�
�
� �f�j�(���ƾ�E9��h_�D���|�_�u�u��o�(�������T��N�U¡�%�d�`�3��l�C���Y����R��1�����'�&�g�3��m�C���P���F��\�����
�b�d�%�w�`�_���&����U�� Y�����'��;�0��1�(�������lW�� 1��\�ߊu�u�
�g��l����I�֓�F�F����
� �d�b��o����+����9��[1�����g�3�
�e�c�-�^�ԜY�Ƽ�T��^1��*��f�%�u�h��0�(�������W��N��ʇ�;�0�
�9��8��������9��UךU���
�`�i�u��>�(�������F��E��AҊ�4�!�'�2�c�m�L�ԜY�����1��*���u�&�<�;�'�2����Y��ƹF��h_�����9�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���Kù��^9��d��Uʷ�2�;�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h_�\���=�;�_�u�w�}�W���Y����l��A��I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�-�Fځ�	����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����lW��G1�����
�<�u�&�>�3�������KǻN��*ۊ�%�#�1�<��4�(�������A	��N�����&�%�d�4��1�[Ϯ�H����E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u����������[��=N��U���u�u�u�
��-��������TF���*���#�1�_�u�w�}�W������F�N��Uʥ�d�4�
�9��3����E�Ƽ�9��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����Z��D��ʥ�:�0�&�u�z�}�WϮ�H����@��V�����'�6�o�%�8�8�Ǯ�H�Ƽ�9��R	����4�
�9�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����R��[
��U���;�_�u�u�w�}�W���&¹��l��R����_�u�u�u�w�1��ԜY���F�N��D���
�<�u�h�'�l����B���F���U���u�u�u�0�3�-����
��ƹF��h\��@���
�g�m�%�w�`�}���Y���R��X ��*���a����w�5����
����A��V�]���h�r�r�u�;�8�}���Y���R��X ��*���a�e�_�u�w�p�W���&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��V�����;�&�2�4�$�:�(�������A	��D��*؊�%�#�1�u����������TOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�g�4�
�;�t�W������F�N��Uʥ�g�4�
�9��3����E�Ƽ�9��h��N���u�u�u�0�$�}�W���Y���F��h\�����1�<�
�<�w�`��������W9��R	�U���u�u�0�1�>�f�}���Y����C��R�����u�%�g�<��)�1���5����@9��h]�G���u�h�_�u�w�}�W���&����Z��_��]���
�e�
� �d�o�(��I���W����ߊu�u�u�u�"��(��@����9l�N�U���
�;�&�2�6�.��������@H�d��Uʥ�g�<�
�<��.����	����	F��X��¥�g�u�
�
�%�:�W���&����_�N�����;�u�u�u�w�4�W���	����@��X	��*���u�
�
�%�!�9�^Ϫ���ƹF�N��U���
�
�;�&�0�a�W���B���F����ߊu�u�u�u�w�}�(݁�����Z�G1�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�'�n�(�������
U��N�U¶�'�,�d�3��m�B���Y����a��R_�����;�&�`�'�0�i�E���s���C9��h�����g�d�%�u�j�u����&����lU��1��U���u�4�2�d�6�1����&Ź��lU��1��\�ߊu�u�
�m�>�;�(��I����[�T�����
�f�e�%�w�3�W�������U��V�����_�u�u�
��(�@���	���l�N��Uʴ�
�:�&�
�!�e�D���?ӑ��]F��D ��*ۊ� �`�g�%��t�J���^�Ʃ�@�N��U���4�
�:�&��+�O��s���C9��h�����e�d�%�u�j�u����K����l	��D1�����a�g�u�;�w�0�(�������P��G�U���%�a�
�g�1��E���	���N��Y	��*���
�;�&�a�1��E���	�ƭ�WF��G1�*���f�`�
�g�l�}�W���YӖ��l��R�����9�2�6�#�4�2�_�������Z��SF��*ڊ�a�
�
�
�8�9����M����U��Uװ���u�x�%�a�2�m�����ƭ�@�������{�x�_�u�w��(���&����_��D�����:�u�u�'�4�.�_�������C9��P1������&�g�
�$��N�ԜY�Ʈ�T��N��U���<�u�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�g�;���P����[��=N��U���u�u�u�
���(������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�
�
�
��-����E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�-�C���H���P
��y*��4���0�8�g�g�2�l����M����9l�N�U���
�
�
�%�!�9�����Ƽ�\��D@��X���u�%�a�0�f�<�(���&����T��E��Oʥ�:�0�&�4��8�W���
����@��d:�����3�8�d�|�w�}�������F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���g�
�&�
�n�t�W������F�N��Uʥ�a�0�d�4��1�W������]��[����_�u�u�u�w�1��ԜY���F�N��A���d�4�
�9�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u����������@��V�����'�6�&�{�z�W�W���&ƹ��l��h�����4�&�2�
�%�>�MϮ�������h�����u�
�
�%�!�9����P�����^ ךU���u�u�3�}�6�����&����P9��
N��@���
�9�|�u�?�3�}���Y���F�G1�����9�
�;�&�0�a�W���&����_��N��U���0�&�u�u�w�}�W���YӖ��l��A�����<�u�h�%�b�<�(���&����l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���%�`�<�
�>�}����Ӗ��P��N����u�
�
�;�$�:��������\������}�
�y�%�b�-���	�ӓ�C9��SGךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�%�`�6�����Y����l�N��U���u�%�`�<��4�W��	����F�N�����u�u�u�u�w�}�WϮ�L����@��S��*ߊ�'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�W���&Ź��F���*���<�
�0�!�%�/����Q����V��C1��A���0�e�$�|�d�t�L�ԶY���F��1��E���
�9�u�&�>�3�������KǻN��*܊�
�
�%�#�3�<����&����\��E�����%�6�y�4��4�(�������@��h��*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C\�����d�|�|�!�2�}�W���Y���F��hX��*ڊ�%�#�1�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����lP��h^�����1�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]ǑN�����0�d�i�u�#�m�C����ד�]ǑN��X���
�
�
�
�'�+�Ͽ�
����C��R��U���u�u�%�c�2�l��������@��h����%�:�0�&�6�����	����l��F1��*���e�3�8�d�~�}�Wϼ���ƹF�N�����}�%�6�;�#�1����H����C9��N�����%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��d�^������F�N��U���%�c�0�d�6�����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����0�d�4�
�;�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�u�w��(���Y����G��X	��*���!�'�'�&�-�u����ۊ��9��1��E���|�f�|�n�]�}�W��Y����V9��V�����&�<�;�%�8�8����T�����h��*���#�1�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����֓�@��GךU���0�<�_�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���!�0�u�u�w�}�W���YӖ��l��h�����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϮ�A����l��A��I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B���F��1��D��u�!�e�a�b�8�F���B���F���*���
�%�#�1�6�.��������@H�d��Uʥ�m�0�d�4��1�(�������A	��N�����&�4�
�0�w�-��������`2��C\�����d�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��Gڊ�&�
�l�|�w�5��ԜY���F�N��M���d�4�
�9�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��1��D���
�9�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���
�0� �!�f���������9��R��]���
�a�
� �e�o�(������C9��Y�����d�n�u�u�'�����&¹��lT��1��U��3�%�-� ����������J9��1�����m�`�%�}�a�9� ���Y���9F������!�g�3�
�d��E��Yۋ��l0��h��C���%�u�;�u�:��Eہ�����l��d��Uʥ��&�9�
��(�F��&���F��S1�����#�6�:�}�2�4�ǫ�
����WN��G1��*��m�%�|�`�~�f�W���	����F
�� 1��*��
�d�i�u�#�����&����\��R�� �&�2�0�}�:��@���&����CU�Z��N���u�%��&�;��(�������S��N�U���
���,�"�����	����R��h��G��
�g�`�u�8�3���P���F��e�����
� �d�c��o�K�������l ��_�*��4�1�!�%�b����Lƹ��]ǻN��*���g�d�
� ��(�E��&���FǻN��U���%�6�;�!�;�l�(ޘ�?�ƻ�V�U�����<�<�
� �e�l�(��I���W����ߊu�u�u�u��<�E��&����R��G]�U���%��9�
�a�;�(��@����[�N��U���%��9�
��(�(���K����CU��_��]���
�8�g�
�"�o�Aہ�K���F�G�����_�u�u�u�w�8�(���Kǹ��lT��1��N���u�%��9��d����A�ӓ� F�d��U���u�!�%�d�n�/���N�ƻ�V�D�����`�'�2�f�g�u�^��^���V
��d��U���u�&�9�!�'�i����A�ѓ� ]ǻN��*���g�d�3�
�c�j����D���F�N��*���&�
�#�a�o�m�G������F��E�����'�2�a�g��t�J���^�Ʃ�@�N��U���%��9�
�g�/���H��ƹF��h8��G��d�8�-�3��l�E���Y���F�N�����:�&�
�#�e�j�1���?�ƻ�V�U�����<�<�
� �d�i�(��I���W����ߊu�u�u�u��<�E��&����R��G\�U���%��9�
�g���������9��R�����u�u�u�%�4�3����J����u ��q(�����}�'�0�2���C���&����l��G��U��|�0�&�u�w�}�W���	����9��h��F��
�g�_�u�w�����K����K9��h\�E���u�h�_�u�w�}�W�������l
��1��3���u�=�;�}�%�8����&�ԓ�F9�� X��G��u�u�d�|�2�.�W���Y�����V��Fڊ�0�
�e�g�]�}�W����ԓ�9��h]�A���u�h�4�
�8�.�(���L����vN��C��U���;�:�e�n�w�}��������l ��\�*��i�u�
�4�e�o�(���J����CT�N�����u�e�n�u�w�-�!���&����l ��_�*��i�u�u�u�w�}��������_��hV�E��e�"�0�u�"�9�����Փ�F9��W��G��u�u�d�|�2�.�W���Y�����V��@ۊ� �f�a�
�e�W�W���&����lT��B1�Bӊ�f�i�u�u�w�}�WϪ�	����U��[�����=�;�}�8�����J����V�
N��R���9�0�_�u�w�}�W���&�ӓ�F9��V��F�ߊu�u�
�4�e�n�(���K����CT�
N�����2�6�#�6�8�u��������l0��1�*���g�l�
�a�w�}��������^��1��*��c�%�|�n�w�}��������T��B1�Aӊ�f�i�u�u�w�}�WϿ�&����G9��\��E��e�e�"�0�w�(��������l ��]�*��e�u�u�d�~�8����Y���F��h8��G���
� �f�e��o�}���Y����_T��h��D��
�g�i�u�#�����&����\��Y�����%��9�
��(�F��&���F��D�����8�
�e�3��i�D���P��ƹF��h8��G��
� �g�l��n�K���Y���F��h8��G��
� �
� �e�e�(��������R�����
�:�
�0��m�N��Y���O��[�����u�u�u�
�6�o�F���&����l��=N��U���4�g�a�
�"�o�G݁�J���9F�N��U����9�
� �e�e�(������	��T��G���
�c�c�%��t�J���^�Ʃ�@�N��U���3�%�;�1��8���O����F9��Y��D�ߊu�u�
�4�e�i����M�ӓ� F�d��U���u�!�%�g��(�F��&����[����*���d�
� �d�`��E��Y���O��[�����u�u�u�0��0�F܁�����9��d��Uʥ��9�
�d�1��G���	�����h�����0�!�'� �$�:����&����lS��E��A��|�~� �&�0�8�_���&�֓�F9��\��D���_�u�u�
�6�o�B܁�����9��R�����9�2�6�#�4�2�_���������V��@؊�0�
�d�f�w�}��������^��1��*��d�%�|�n�w�}��������l ��]�*��i�u�u�u�w�}��������9��O1��*��d�%�u�=�9�u��������9��C1��*��`�%�}�|�j�z�P������F�N�����9�
�
�g�1��D���	��ƹF��h8��G���d�
� �g�d��D��Y���F� ��&���
� �g�g��n� ���Yۉ��P	��1��*��c�%�}�|�j�z�P������F�N�����0�a�3�
�`�j���Y����l0��1�����g�f�%�u�j�W�W���Y�ƭ�l��D�����e�"�0�u�#�-�F������� N��S��D���0�&�u�u�w�}�WϿ�&����G9��Z��E��e�_�u�u��<�E�������F9��X��F��u�u�u�u�w�<�(���
����R��q(��3ʢ�0�u�7�8�%�8��������
T��F�U���d�|�0�&�w�}�W���YӖ��R
��1����`�n�u�u�'��݁�&����V��G\��Hʦ�1�9�2�6�!�>��������V��h8��G���'�2�f�b�~�v��������G��Y�� ��l�
�d�|�]�}�W����ԓ�l ��Y�*��i�u�u�u�w�}��������G��h[�*��� �g�`�
�f�*��������]��B1�Bي�g�e�u�u�f�t����Y���F� ��&���3�
�c�b�'�f�W���	����9��Q��B���%�u�h�_�w�}�W�������9��h\�A���u�=�;�}�%�>��������
P��F�U���d�|�0�&�w�}�W���Yӈ��`��h��G���
�f�_�u�w�����@����S��G]��H�ߊu�u�u�u�:��Fׁ�����l��@��U¡�%�a�
� �`�o����P���A�R��U���u�u�u�%�d�;�(��&����F�G1��؊�
�d�3�
�f�e����D���F�N��#���
�e�
� ��(�D��&����[�������:�
�
�:��(�D��&���F�_��U���0�_�u�u�w�}�(���K�ԓ�9��h]�E���n�u�u�%��1�(�������9��R�����u�u�u�%�4�3����H˹��D��F����
�0�
�m�d�m�W���H����_��=N��U���u�%�6�;�#�1�Fׁ�I����9F���9���
�:�
�:�'�>��������9��R�����9�2�6�#�4�2�_�������]��Y�����
�!��'��2�(�������9��B�\��u�u�%�<��)�1���5����@9��h]�E���u�h�_�u�w�}�W�������l
��1����u�!�%�d�e�;�(��K����O�I�\ʰ�&�u�u�u�w�}����H�֓�F9��W��D�ߊu�u�
�:��l����I�ޓ�F�F�����1�/�'�&�d�;�(��I����K	��V�����
�#�
�|�]�}�W�������l ��\�*��i�u�1�9�#�9����
�ғ�F9��Z��Fʭ�'�4�
�:�$��ށ�P���F��Y�����
�a�c�%�w�`�_�������I��D1�����f�m�%�u�8�}��������EW��UךU���
�%�
� �o�o����Dӕ��l
��^�����'�&�2�0��-��������lU��C�����1�!�%�d�f�;�(��&���l�N����� �d�f�
�e�a�W���&����P9��T��]���;�1�4�
�8�.�(���&���F��P ��]���
�a�3�
�d�n����B�����h��G��
�f�i�u�w�}�W�������]��[��Dʢ�0�u�!�%�o�����I���F�_��U���0�_�u�u�w�}��������EU��d��U���u�%�&�
��<����&����CW�
N�����2�6�#�6�8�u����ە��]��G��*ۊ� �l�a�%�~�n�^��s���C	��h_�� ��a�%�u�h�$�9��������G	��B �����}�%�6�;�#�1�F݁�P����]��Y��3؊�
� �c�c�'�t�L���Y�����1����� �d�d�
�f�a�W���&����P9��T��]���<�0�&�2�2�u��������W��G�G���_�u�u�%�$����H¹��Z�D�����6�#�6�:��3����ۇ��P	��C1��D؊�|�~� �&�0�8�_�������U��UךU���u�u�:�g�f�>��������l��S�����:�<�
�0�#�/�����ο�T����G���3�
�`�
�e�q�E���s�����1�����`�
�g�i�w�)�(�������P�������1�4�
�:�$�����J���F��P ��]���d�3�
�`��o�^�ԜY���F��D\�����3�
�`�`�'�}�Jϭ�����Z��R��§�&�/�}�<�9�9����&����T��G\��F���n�_�u�u�8�o����L�֓�F���*���<�
�0�!�%�(�����έ�l��D�����f�u�u�;�>�3�ǘ�&���� ^��G�U���$�
�
� �`�o����D���F�N�����d�3�
�l��n� ���Yے��lS��Q��@Ҋ�g�e�u�u�f�t����Y���F���*��
� �b�a�'�f�W�������@��h_�� ��l�
�g�i�w�/��������
W��N��ʤ�
� �d�d��n�L���Yӗ��R��P ��*���d�l�
�g�k�}����¹��T9��\�����7�d�'�2�d�e�^�ԜY�ƽ�l��^	��@���
�f�e�%�w�`�_���&�ԓ�F9��Z��Gʴ�1�$�<�
�"�o�Gہ�J��ƹF��U1�����
�
� �f�d��E��Y۔��l��Q��E���%�u�;�u�5�)�F�������O��N�����&�<�;�l�1��F���	���N��^1��*���f�l�
�g�6�9����&����T9��V����u�7�3�
�d�m����D���F�N�����'�2�f�e�w�5��������l ��\�*��e�u�u�d�~�8����Y���F��Z��M���
�f�g�%�l�}�Wϯ�����lT��1��U��%��9�
�`�;�(��M����
F��@ ��U���_�u�u�
��(�O���	���N��G1�*���b�e�%�u�9�}����O����R��G\����u�
�
� �e�l�(��E���F��R �����d�l�3�
�d�l����Y����\��h��*���0�&�u�d�l�}�WϬ�J���� V��h�I���e�u�=�;��0�(��&����W��S�����;�!�9�g��t����Y���9F���*���f�m�
�g�k�}�G������G��[�����a�`�u�u�'�>��������O��[��W���_�u�u�
�����MŹ��Z�D�����6�#�6�:��5��������F��P ��]���6�;�!�9�b��1���?����u ��B��*���0�0�}�;�>�3����^����^��1��*��c�%�}�d�f�9� ���Y���O��N�����a�3�
�m�o�-�W��
����\��h�����&�2�0�}�:��C���&����l��E�����1�!�%�m��(�E��&���l�N��#���3�
�m�g�'�}�Jϭ�����Z��R��¦�2�0�}�8��k����A�ޓ�O������!�%�m�
�"�o�Eہ�H����F�E1�����c�l�%�u�j�.��������V��EF�����'�2�!� �$�:����	����@��A[��F��������t��������AN��D�����e�u�u�8��d����O�ߓ�N��_�����:�e�|�|�l�}�WϬ�����U��N�U¡�%�d�
� �f�l�(������^��1��*��b�%�|�_�w�}�(���H����P��G\��H���8�
�g�
�"�e�E���Y����lW��B1�M���|�_�u�u���E���&����l��S�����d�d�3�
�d�j����Ӕ��l ��]�*��n�u�u�'�>�4�(���J����CT�
N�����a�
�0�
�f�m����&����lU�� 1��\�ߊu�u�
�
�c�;�(��H����[�C��D���'�2�a�c�w�/��������P��G�U���'�<�<�3��n�F���Y���G��]�� ��m�
�d�:�w����N����]ǻN�����3�
�`�d�'�}�J�������9��h_�F���u�:�u�%�4�3����H���9F���G���
�b�
�g�k�}����H�ԓ�F9��1��U���u�%�6�;�#�1�F��B�����1��*��m�%�u�h��0�(��&����W��G]�����%�6�;�!�;�l�F��Y����V��Q��@���%�u�h�}�8�1����6����A��R����� �9�&�3��h�G���Y����R��X ��*���
�|�_�u�w�8�O���&����l��S�����d�l�'�2�d�d�W���Y����\��h��*���_�u�u�0�n�;�(��O����[�C��D���3�
�c�m�'�}����	����@��A_��\�ߊu�u�0�
�"�l�Bށ�K�����hV�����`�f�%�u�8�}��������EW��UךU���0�
�8�d��(�F��&���FǻN��U���
�4�g�f�1��C���	�ƻ�V�D�����
� �d�a��o�G���Y�����RNךU���u�u�0�
�:�j����M�ד� ]ǻN�����8�d�
� �f�h�(��E����^��1��*��l�%�u�:�w�-��������lW�=N��U���
�8�d�
�"�l�A߁�K�����h��L���
�a�`�%�w�3�W���&����9��h_�A���|�_�u�u�2����L����\��Y1��*��`�%�u�h��0�(�������P��X�����
�0�
�l�b�f�W���
����^��h��D��
�f�i�u�w�}�W���	����9��Q��A���%�u�=�;��8�(���H����lW��1��]���h�r�r�u�;�8�}���Y���@��C��E���
�a�c�%�l�}�Wϭ�����R��B1�Bފ�g�i�u�d�w�5�������� ��E��F��|�i�&�2�2�u��������EW��X��U���0�w�w�_�w�}��������l��X�����
�c�c�%�w�`�_���	����lT��1��U���'�#�
� �e�j�(��B�����h��D���1�8�'�4��(�E��&���F��R����d�1�8�'�6����IŹ��	��C��Bӊ� �g�b�
�e�f�W���
����^��h��D��
�g�i�u�$�1����M����R��h����!�%�&�3��o�O���P���F��[1�����3�
�c�f�'�}�J�������l ��[�*��:�u�8�
�n�3����&����l��d��Uʦ�9�!�%�b�1��A���	���N��G1�*���d�c�
�g�6�9��������l ��X�*��n�u�u�&�;�)��������S��N�U���u�u�u��9�8�(���&����lW��B1�B݊�g�"�0�u�$�1����N����P��h�E���u�d�|�0�$�}�W���Y����V��B1�@ۊ�g�_�u�u�2����&����T��G]��H�ߊu�u�u�u�6�:�F�������\��B1�@݊�g�"�0�u�$�1����N����P��h�E���u�d�|�0�$�}�W���Y����lW��h�� ��m�
�g�_�w�}�����ד�F9�� Z��F��u�u�u�u�w�-��������l*��G1����� �f�`�
�f�*����
����^��B1�Cӊ�g�e�u�u�f�t����Y���F���*���9�
�:�
�8�-����&����l��=N��U���
�8�g�
�"�o�Fف�K�����h\�����f�b�u�:�w�-��������lW�=N��U���
�8�g�
�"�o�Dށ�K�����1��*��c�%�u�;�w�.��������^�=N��U���
�8�g�
�"�o�Dف�K�����h\�����f�b�u�;�w�.��������^�=N��U���
�8�g�l�3�0����&����U��G\��H���8�
�l�3��n�O���Y����^��^�� ��e�
�g�n�w�}��������l ��\�*��i�u�u�u�w�}��������U��\�����=�;�}�8��o����K�֓�N��S��D���0�&�u�u�w�}�WϮ�/����9��P1�@��u�u�&�9�#�-�Cف�����R��B1�AҊ�g�i�u�&�;�)���&����A��h��F��
�g�:�u�:��Gށ�����9��UךU���0�
�8�g��(�E��&���FǻN��U���0�
�8�g��(�E��&����[����*���c�
�0�:�0�3����K�ԓ�N��S��D���0�&�u�u�w�}�WϮ�/����9��P1�@��u�u�&�9�#�-�B���&����l��S�����d�'�2�f�e�}����	����@��A_��\�ߊu�u�0�
�:�o�(���K����CT�
N�����3�
�g�m�'�}��������V��[�N���u�&�9�!�'�j����N����Z�=N��U���u�8�
�d��(�A���	�ƻ�V�C��Aۊ� �c�g�%��t�J���^�Ʃ�@�N��U���4�
�:�&��+�O��s���@��C��M���
�m�
�g�k�}����M¹��lP��h����4�
�:�&��+�(���s���@��C��L���
�m�
�g�k�}�&���&����9��hX�*��4�1�&�9�#�-�O���&����CT�=N��U���
�8�g�3��k�E���Y���G��^�����c�f�%�u�8�}��������EW��UךU���0�
�8�f��(�F��&���F��R����
�0�
�l�e�<�Ϫ�	����l��h]�C��u�u�&�9�#�-�G�������Q��h�I���&�9�!�%��(�F��&����\��G1�����9�d�d�n�w�}��������l ��V�*��i�u�u�u�w�}��������U��^�����=�;�}�0��0�D߁�����9��^��H��r�u�9�0�]�}�W���Y����G�� 1����l�n�u�u�$�1����K����^��h�I���!�%�d�c�%�:�D��Y����R��X ��*���
�|�_�u�w�8�(���J����lW��1��U��}�0�
�8�e�����@����]��R����
� �d�g��o�L���Yӕ��l��Z�� ��f�
�f�i�w�}�W���YӖ��R
��1��*��f�%�u�=�9�u��������U��]�����|�h�r�r�w�1��ԜY���F��[1�����3�
�m�e�'�f�W���
����^��h��L���%�u�h�}�4�-�(���@�ԓ�F��SN����
� �b�m�'�t�}���Y����G��1��*��e�%�u�h��0�(��&����V��N��U���
�b�;�!�1��F���	����F�D�����b�3�
�d�a�-�W��Q����^��B1�L܊�g�4�1�&�;�)��������V��G�U���&�9�!�%�o�;�(��K����[�N��U����;�0�
�;�����J����V��h����u�&�9�!�'�j����H�Г�N��S��D���0�&�u�u�w�}�WϬ�����l_��h����u�0�
�8�d����M˹��Z�=N��U���u�4�2�d�6�1����
�ԓ�F9��Z��Gʢ�0�u�&�9�#�-�@���&����l��G��U��|�0�&�u�w�}�W���	����l��Q��D���%�n�u�u�$�1����&����^��G\��H���0�m�'�2�c�l�W���Y����G��h��F��
�g�n�u�w�.����	�֓�F9��]��G��u�!�%�`��8�(��HӞ����T�����d�d�n�u�w�.����	�ד�F9��^��G��u�!�%�e�1��N���	�ƭ�WF��Y��D���2�f�`�|�]�}�W���&����9��h_�@���u�h�}�8��d����J����R��^�����'�2�f�`�~�W�W�������CR��Q��E���%�u�h�_�w�}�W���&����l��B1�Aߊ�f�"�0�u�#�-�@߁�����9��^��H��r�u�9�0�]�}�W���Y����_T��1��*��`�%�n�u�w�.����	�ғ�F9��W��F��u�u�u�u�w�.����	�Փ�F9��Y��Fʢ�0�u�&�9�#�-�Dځ�����R��B1�Cߊ�g�e�u�u�f�t����Y���F������d�
� �d�c��D�ԜY�ƿ�_9��GZ�����e�b�%�u�j�u����A����lU��N��ʴ�
�:�&�
�!��^�ԜY�ƿ�_9��GZ�����e�m�%�u�j�u���&����^��G\�����6�%�
�0��d�B��Y����V
��Z�*���g�l�
�g�k�}����J����S��h����4�
�:�&��+�(���s���@��C��M���
�c�e�%�w�`�_���N����S��h����&�9�!�%�`�;�(��M����l�N�����%�l�3�
�a�e����D�ή�\
��p+�� ���'�4�0�
�%�����
����S��h����<�8�f�
�8����H����]ǻN�����8�a�3�
�a�n����D���F�N��G���
�<�u�=�9�u�����Փ�F9��V��G��u�u�d�|�2�.�W���Y�����h��D���
�c�a�%�l�}�Wϭ�����V��B1�Gފ�g�i�u�!�'�j�(���K����CT��Y
�����8�a�
� �e�l�(��B�����h��@ۊ� �g�f�
�e�a�Wǭ�����S��S�����
� �g�f��o��������]��[��D��u�u�&�9�#�-�E���&����l��S�����m�
� �g�o��EϿ�ӕ��l��_�� ��f�
�g�n�w�}��������l ��Y�*��i�u�u�u�w�}��������_��N�����&�9�!�%�o�/���L����[�I�����u�u�u�u�w�<�(���
���� 9��=N��U���
�8�`�
�"�o�O؁�J���9F�N��U���
�8�`�
�"�o�O߁�Jӑ��]F��E1�����3�
�c�a�'�u�^��^���V
��d��U���u�%�&�3��k�A���B�����h��@ߊ� �g�l�
�d�a�W���Y�����T�����f�f�"�0�w�.����	�ԓ�V��X�E���u�d�|�0�$�}�W���Y����C9��Y�����c�_�u�u�2����&����W��G\��H���8�
�l�3��n�O���Y����R��X ��*���
�|�_�u�w�8�(���LĹ��lU��1��U��}�8�
�e��(�D��&����]��R�����
� �f�d��o�L���Yӕ��l��V�� ��f�
�g�i�w�.����	����W��E	��*���f�f�
�g�/�/��������_��G�U���&�9�!�%�n�;�(��K����[�C��D���3�
�a�m�'�}��������CS��Q��A���%�|�_�u�w�8�(���L����R��h�I���&�9�!�%��(�F��&����]��Z��D���
�f�l�%�~�W�W�������CP��Q��A���%�u�h�}�2����O����\��Y1��*��m�%�u�:�w�-��������lW�=N��U���
�8�c�
�"�n�A߁�K�����h_�*���f�d�
�g�6�9��������l ��Z�*��n�u�u�&�;�)��������T��Q��G���%�u�h�}�:��(���&����	��^��*���
�m�e�n�w�}��������U�� ^�����h�}�8�
�b�����N����]��R�����c�c�%�|�]�}�W���&����l ��Z�*��i�u�u�u�w�}����Hʹ��lW��1��U���;�}�8�
��(�F��&���F�_��U���0�_�u�u�w�}��������ET��UךU���0�
�8�m�1��C���	���N��G1�����g�f�%�u�8�}��������EW��UךU���0�
�8�l��2�(���H����CT�
N�����8�f�
� �f�l�(������C9��Y�����d�n�u�u�$�1����&����U��G\��H��� ����%�:�D��Y����@��C��*���d�g�
�g�l�}�Wϭ�����l ��X�*��i�u�!�%�f�h����O�Փ�F��SN��Ҋ�0�
�g�d�l�}�W���Yӕ��R��1����� �c�m�%�w�`��������l��C�����/�}�<�;�3�.�(���&¹��lP��h�Y��|�_�u�u�$�����&����V��N�U���u�u�u�!�'�n�(���O�ޓ�F��R ��$���
��
�
�"�k�E���Q���A��N�����u�u�u�u�#�-�C߁�����l��=N��U���u�=�4�!�4�.�(���H����CW�
N�����2�6�#�6�8�u����ە��]��D����� �d�d�
�d�q�E���s�����V�����g�g�%�u�j�W�W���Y�Ƹ�C9��Q��G���%�u�=�;���9���:����lU��F�U���d�|�0�&�w�}�W���YӒ��lS��B1�E݊�g�_�u�u�>�3��������U��[�����h�_�u�u�w�}����@����_��h����u�&�9�!�'�o����@�ӓ�N��S��D���0�&�u�u�w�}�Wϭ�����W��B1�@ڊ�g�_�u�u�>�3��������]	��Q��E���%�u�h�}�>�3��������U��[�����:�u�%�6�9�)����H��ƹF��^	�����2�
� �g�c��D��Y���F���*���3�
�d�e�'�}����Q����G��1��*��c�%�}�|�j�z�P������F�N�����!�%�d�3��l�F���B�����Y1�����
�:�
� �e�d�(��E����Z��V����� �g�a�
�d�%�Ͽ�&����G9��1�N���u�&�2�7�#�;�(��A����[��h8��G��
� �f�`��o�D�������U��d��Uʡ�%�e�3�
�n�i����D�΢�D��Y��*ۊ� �d�c�
�d�<�ϭ�����V��B1�Fي�g�n�u�u�#�-�F���&����l��S�����3�:�
�
�"�l�Oց�KӉ��@��h�����d�;�!�3��m�N���P���F��G_�����e�g�%�u�j�u�����ד�F9��_��Gʴ�1�&�9�!�'�h����I�ѓ�O��N�����f�3�
�a�e�-�W��Q����Z��^��*���g�`�
�f�8�}����O����U��h�N���u�!�%�a�1��F���	���N��G\�*���:�2�;�3��l�@���Y����R��X ��*���
�|�_�u�w�0�Fځ�����9��R��]���0�2�a�
�2�2����¹��lU��1��U���!�%�l�
�"�n�F߁�K��ƹF��Z�*���f�d�
�g�k�}����@ʹ��^	��V �� ��e�
�g�-�%�<�(���
����9��d��Uʡ�%�b�3�
�d�d����D�ή�^��RZ�����'�4�
�g�1��D���	�ƣ���hW�����g�l�%�|�]�}�W���H˹��lU��1��U��&�1�9�2�4�+����Q����T����*���&�2�u�u�9�4����	����9��h��*��e�|�_�u�w�0�F���&����l��S�����m�
�0�:�0�3����M�Փ�F��EN��*���&�
�#�
�~�W�W�������l��X�����
�a�f�%�w�`�_���&�Г�F9��]��Fʺ�u�0�
�8�f����Nʹ��]ǻN����g�6�&�
�6�)����Lǹ��Z�=N��U���u�%�6�;�#�1�F݁�Y����N��v ��;��� �`�m�%��t�J���^�Ʃ�@�N��U���4�
�:�&��+�E��s���G��V�����2�;�3�
�o�l����D�θ�C9��1��*��m�%�u�'�$�1����L����lU��G�U���!�%�m�
�6�)����&����R��N�U���u�u�u�4��2�����ԓ���YN�� �����d�3��k�(��I���W����ߊu�u�u�u�'�>��������]ǻN����`�1�8�'�6����Jù��Z���M���3�
�a�e�'�}�ϼ�����V��R�����<�3�
�a�c�-�^�ԜY�Ƹ�CT��h
�����;�3�
�d�`�-�W��Q����l��Q��E���%�u�'�7�:�/��������T��^_�� ��g�
�g�n�w�}����@ʹ��^	��V �� ��e�
�g�i�w�-�Dׁ�K���� T��h����'�0�2�a��8��������U��^�����_�u�u�8�e�;�(��H����[�[*�� ��c�
�d�4�3�/����&����l��d��Uʡ�%�
� �d�c��E��Yە��l��[�� ��b�
�g�:�w�8�(���Jù��G9��h_�B���|�_�u�u�:�i����H�Г�F�F�����;�<�
�0��d�DϿ�ӕ��l��^�� ��d�
�g�n�w�}����&����V��G\��H���#�'�9�"�1��F���	�ƣ���Y1�����
�:�
� �e�d�(��B�����1��*��m�%�u�h��/����&����W��G\�����0�
�8�g��(�E��&���9F���B���
�m�c�%�w�`�_���K�ޓ�V��P�����m�d�%�u�8�}��������EW��UךU���8�m�3�
�n��E��Yۊ��9��hW�*��4�1�'�#��(�N���	����F�C��*���d�m�
�g�k�}��������l��h]�Mʺ�u�0�
�8�n���������9��UךU���8�
�e�
�"�n�G܁�K���W�@��U �
�&��&��)��������9��P1�B���u�%�6�;�#�1�D��Y����D��d��Uʡ�%�d�d�3��i�O���Y���D��_��]���6�
�4�0��/��������l��hZ�@��4�
�:�&��+�(�������V�=N��U���
�e�
� �d�l�(��E���F��R �� ���&��&�
�#�(����&����A��^�U���%�6�;�!�;�n�A������D��N�����d�a�3�
�a�i����Dӕ��l
��^�����'�'�&�/��3����ۏ��_��X�����&�'�2�a�n�q�C���s���G��^�����c�f�%�u�j��Uϩ�����Z��SF�����d�a�
�e�w�}����ۖ��l��D��\ʰ�&�u�e�n�w�}����H�Г�F9��V��A��u��-� �.�(�(��&����W��G\��Dʱ�"�!�u�|�]�}�W���Y����V��B1�Cߊ�d�i�u�!��2����������^�����0�}�8�
�n�;�(��A����U��UװU���!�%�d�e�1��B���	�����1��*���e�%�}�d�3�*����H��ƹF��Z��Dۊ� �d�b�
�d�a�W���H����S��h�D���:�;�:�d�~�W�W�������9��h[�*��i�u�'�2��l����Aǹ��P��N����!�u�|�_�w�}����HŹ��lP��h�I���'�2��d�1��Oہ�H����F��S�����|�_�u�u�:��F؁�����l��S�����
�
� �c�e�-�_��T����\��XN�N���u�!�%�d�o�;�(��&���F��G1�*���b�m�%�}�o�p�FϺ�����O��N�����d�l�3�
�c��F��Y����_��B1�E���}�m�x�d�3�*����P���F��G1�*���d�c�
�g�k�}��������E��X�����
�0�!� �$�:��������l ��\�*��y�:�<�!�0�/��������V�N��*���
�4�!�3��o�N���Q�����Y��E���|�n�u�u�#�-�F�������9��R������c�3�
�c��DǪ�&����T��B �����}�8�
�c�4�.�(���N�֓�O�S�����:�<�!�2�%�(�����θ�C9��h�����
�b�
�d�~�}����Q����]��R�����;�1�!�%�a���������9��G�U���;�u�:�<�#�:�ǫ�
����WN��G1�*���!�3�
�b��l�^��J�Ʃ�@�L�U���!�%�d�d�1��Gׁ�H���G��Z�� ��c�%�}�u�w�}�������9F���*��
� �m�m�'�}�J�ԜY���F��h�����#�
�u�=�9�u����L����V��G\��\��r�r�u�9�2�W�W���Y�Ƽ�\��Q��D؊�g�_�u�u�:��E܁�����l��S�����:�<�
�0�#�/�����ι�@��R
�����g�
� �m�o�-�^��P��ƹF��Z��Gފ� �m�e�%�w�`��������l��C�����!�'�2�!�"�.����Q����\��h��A���������^ê�&����T��B �����}�e�u�u�:��E܁�����l��_��U���;�:�e�|�~�f�W�������Q��B1�G���u�h�%��;��(���N�֓� N��N����!�u�|�_�w�}����K˹��lW��1��U��%��9�
��(�F��&���F��@ ��U��n�u�u�!�'�l�N���&����CR�
N��*ۊ� �c�c�%��l��������l�N����
� �d�m��o�K���H�ƻ�V�D�����8�
�
� �f�m�(��Y�ƿ�T�������!�9�d�
�a�t����Y���9F���*��
� �l�m�'�}�JϪ�	����U��\��G��u�:�;�:�f�f�W������� T��B1�E���u�h�%�&�����M����W��X����|�_�u�u�:��Dہ�����9��R�����
�
� �l�c�-�_������\F��UךU���8�
�f�
�"�l�Aہ�J���C	��h_�� ��a�%�}�d�3�*����H��ƹF��Z��Fӊ� �g�d�
�f�a�W����ԓ�9��h]�A���}�u�u�u�8�3���B�����h_�����f�
�d�i�w�/��������9��[�X��1�"�!�u�~�W�W�������9��h\�E���u�h�%��;��@���&����l��]�����:�f�|�_�w�}����M¹��lT�� 1��U��%��9�
�`�;�(��M����V��X����|�_�u�u�:��C܁�����9��R�����9�
�d�3��i�D���Q����\��XN�\�ߊu�u�8�
�c����LŹ��Z��������!��2�)����&����_9��Q��@���%�u�u�:�;�%�2ߑ�����R��h!��0���9�d�3�
�b�e����s���G��Z�����m�b�%�u�j�;����,����F��B�����d�a��3��e�B���Q���W��X����n�u�u�!�'�l�(���H����CT�
N�����2�6�#�6�8�u����ۇ��P	��C1��D؊��|�~�&�0�8�_�������U��UךU���8�
�`�
�"�o�@ց�H���U��O#��!���!��9�<�;��E؁�&����S��G\��D���d�1�"�!�w�t�}���Y����S��B1�D݊�g�i�u�d�w�5�������� ��E��F��|�k�&�2�2�u��������EW��Y��U���0�w�w�_�w�}����Où��lU��1��U��7�3�e�d�c��G��Y����W	��C��\�ߊu�u�8�
�a����K˹��Z�U��E��a�
�e�f�w�2����J����F�C��D���3�
�c�g�'�}�Jϼ��֓�R��F^��Dʱ�"�!�u�d�l�}�WϪ�	����U��\�����h�&�1�9�0�>�����ο�T�������!�9�d�
��t�\ϭ�����uT��R	��M��|�_�u�u�:��@���&����l��S��D���=�;�}�<�9�9����HŹ��lW��1��\��&�2�0�}�'�>�������� S������w�_�u�u�w�}����A����G9��h_�M���u�h�&�1�;�:��������A��M�����1�!�%�d��(�F��&��� T�dךU���8�
�m�3��n�@���Y���D��_��]���0� �!�&�1��D���	���R��X ��*���a�e�u�9�2��U�ԜY�Ƹ�C9��h��D��
�d�i�u�6��(���H����CU�N�Dʱ�"�!�u�|�]�}�W���&¹��lS��h�I���d�u�=�;��0�(ׁ�����l��
N��*���&�
�#�f�g�}����[����F�C��Gڊ� �d�e�
�f�a�W���&����P9��T��]���<�0� �&�0�8�_�������]9��Q��F���%�|�g�|�l�}�WϪ�	����U��\��G��u�!�
�:�>�����ۓ��Z��SF����
�4�!�6�$����M����M��Y�����0�%��3��o�(��P���F��G1�*���d�f�
�g�k�}�F������@��R
�����3�
�`�d�'�t�Kϭ�����R��X ��*���g�f�|�u�;�8�U���s���G��]�� ��`�
�d�i�w�0�(ہ�����9��\�X��1�"�!�u�~�W�W�������l ��[�*��i�u�!�
�8�4�(�������V��RF�����0�}�:�d�4�.�(���H����CW�Z��N���u�!�%�g��(�F��&���F��G1�*���d�c�
�g�e�}�W�������V�=N��U���
�c�3�
�b�l����Dӕ��l
��^�����'�&�<�!�%�:�ǭ�����^��a1��*��`�%�|�!��3����Q����T��I�U���8�
�a�3��h�@���Q�����Y��E���|�n�u�u�#�-�E؁�����9��R��W���"�0�u�&�0�8�_���K����S��h�U���<�;�1�4��2�����ԓ�O�R��U��n�u�u�!�'�o�(���H����CU�
N�����3�
�d�`�'�u����������^	��¡�%�d�
�4�#�;�(��A����F��@ ��U���<�!�2�'�"�.����Q����^��V�����g�m�%�|�~�*��������G��EF�����0�}�8�
�o�>��������9��G�U���;�u�:�<�#�:�ǫ�
����WN��G1�*���!�3�
�g�o�-�^��L����_��C�����u�8�
�l�1��A���	�����h�����0�!�'�'�$�'�_���������1����� �d�g�
�f�q�C���s���G��W����� �d�m�
�e�a�WǪ�	����U��W�����:�u�%�6�9�)����H��ƹF��Z��*���d�a�
�d�k�}��������E��X�����0� �&�2�2�u��������G9��h_�L���|�`�|�n�w�}����Jù��lW��1��U��w�w�"�0�w�����&����U��_�����u�%�6�;�#�1�Bہ�PӃ��VF�UךU���8�
�d�3��k�N���Y���D��_��]���g�3�
�`�g�-�W���	����@��A_��F���0�&�u�e�l�}�WϪ�	����U��]�����h�}�8�
��8�(��JӉ��F��E�����
�d�c�%�~�W�W�������l ��_�*��i�u��;�2���������l��1��*��c�%�u�:�w�-��������lW�=N��U���
�a�3�
�d�n����DӒ��lW��Q��F���%�}�u�u�w�2����I��ƹF��Z��@���
�d�a�%�w�`�_�������T9��V�����%�6�;�!�;�l�F��Y����^��1��*��
�d�i�u�#�����&����\��R�� �&�2�0�}�/�����&¹��lP��h�Y��|�_�u�u�:��@���&����CU�
N�����;�!�9�d�f�{����H�Г�F9��1��\�ߊu�u�8�
�o�;�(��&���F�N�����!�%�d�a�1��Oׁ�H����C9��Y����
�|�0�&�w�m�L���YӒ��lU��Q��CҊ�g�i�u�!��2����������Y�����:�&�
�#�e��G���Y����V��1�����`�
�g�|�]�}�W���&����lW��1��U��&�1�9�2�4�+����Q����V��G1�����9�d�
��~�v�����Ί�l��h]�D���_�u�u�8��m����Nǹ��Z�D�����6�#�6�:��3����ۇ��P	��C1��D؊�e�u�u�;�>�3�ǘ�&¹��lP��h�\�ߊu�u�8�
�f�;�(��&���F�N������
�
� �a�k����Y����\��h��G��|�0�&�u�g�f�W�������9��hY�*��i�u�d�u�?�3�_���������V��D���
�m�
�f�w�}��������C9��Y����
�c�|�0�$�}�G��Y����^��1��*��f�%�u�h�]�}�W���Y����\��h��*���=�;�}�8��j����J�ѓ�N��S��D���0�&�u�u�w�}�WϮ�����lW�� 1��N���u�!�%�a��(�@���	���D�������;�<�;�1�$�����&����V��G��U���<�;�1�4��2�����ԓ�O�R��U��n�u�u�!�'�i�(���N�ғ�F���*���<�
�0�!�%�/����Q����T�������d�6�&�
�"�k�O���P����]ǻN�����c�3�
�d��o�K�������T��A�����=�3�
�<�?�u����ۋ��l0��h��C���%�|�!�
�9�8��������V�I��U���
�`�3�
�f��F��T�ƨ�D��^��\���_�u�u�u�w�0�(�������9��R�����9�2�6�#�4�2�_�������Z��SF����b�3�
�l��l�[��P��ƹF��Z��M���
�f�d�%�w�`��������l��C�����/�}�;�<�9�9����M����lW��1��\���|�n�u�u�#�-�Cց�����l��S�����:�<�
�0�#�/��������GN��D�����8�
�b�3��n�(��U����]��R�����;�1�r�r�q�.�(���&¹��@��B1�M���}�d�d�1� �)�W���P����F�C��A���
�g�m�%�w�`��������l��C�����!�'�2�!�$�:��������U��W�����!�
�;�0�2�u�������A���*؊� �d�a�
�f�n�Z�������V�G����u�8�
�e�1��Bׁ�K���W�@��U¦�2�0�}�8��d����O˹��F�D�����%�6�;�!�;�l�(��PӃ��VF�UךU���8�
�d�3��n�B���Y����G��X	��*���!�'�&�<�#�/��������]��V�����
�#�a�f���1���?������^ ����� �&�2�0��m�W�������l ��]�*��f�x�u�:�9�2�G���P��ƹF��Z��G���
�c�
�g�k�}��������E��X�����1�4�
�:�$�����?���F��P ��]���d�3�
�`��o�^�ԜY�Ƹ�C9��h��B���%�u�h�w�u�*����
����WN��h_�� ��c�%�|�k�$�:����	����@��A_��D���u�9�0�w�u�W�W�������l �� W�����h�&�1�9�0�>�����ο�T�������!�9�d�
��t�\ϭ�����uT��h��C���%�|�n�u�w�)���&����T��N�U��u�=�;�}�>�3�Ǫ�	����U��X��G���u�<�;�1�6�����&����lU��N�����e�n�u�u�#�-�Bف�����l��S��E���=�;�}�
�2�(��������9��S�����;�!�9�`��t����Y���9F���*���3�
�b�l�'�}�Jϭ�����Z��R��§�&�/�}�;�>�3�ǯ�&����T��h��D��
�g�y�m�~�W�W�������l ��\�����h�&�1�9�0�>�����ι�@��R
����l�6�&�
�6�)����Hǹ��F�B �����}�-�
�
��(�A���	���9F���*���3�
�c�
�e�a�W��Y����N��P ��]���d�d�3�
�c��E���Y����V��G1�����9�d�
�c�~�8����I��ƹF��Z��*���d�e�
�g�k�}��������E��X�����;�1�4�
�8�.�(���K����K��Y������
�0�
�o�l�^�ԜY�Ƹ�C9��h��L���%�u�h�&�3�1��������AN��D��]���<�;�1�%�$��(�������
S��G_��@���n�u�u�!�'�k�(���H����CU�
N��#���
�
� �d�`��D��Y����G	�G�U���!�%�c�
�"�d�O���Y����G��X	��*���!�'�&�<�#�/����
����WN��Y1��C���
�a�
�f�{�2��������]��Y��R��s�!�%�c��(�N���	����W��X����|�|�n�u�w�)���&���� ^��G_��Hʥ��9�
�
�"�l�@ց�J���W��X����n�u�u�!�'�k�(���H����CT�
N��Wʢ�0�u�&�2�2�u����H����
S��G\��Iʦ�2�0�}�%�4�3����H����O��[��W���_�u�u�8��h����I�Г�F���*���<�
�0�!�%�/����Q����T����G���6�&�
� �n�m����L���9F�N��U���
�c�6�&��(�@���	�����h�����0�!�'�'�$�'�_�������^��1��*��
�g�y�g�~�W�W�������9��h_�F���u�h�%��;��(���H����CT�N�����u�f�n�u�w�)���&����Q��G\��H���w�"�0�u��3�݁�&����lW��1��U���%�6�;�!�;�h�(�������V�=N��U���
�b�;�!�1��F���	���N��G1�*���d�g�
�g�/�/��������_��G�U���!�%�c�
�"�l�Nف�K���W�@��U¥�&�
�
� �n�i����Y����\��h��G��|�0�&�u�g�f�W�������
9��h_�B���u�h�}�4�0�l��������9��h_�����l�g�%�u�8�}��������EW��UךU���8�
�
� �b�o����Dӕ��l
��^�����'�'�&�/��3����ۃ��l��h8�� ���g�%�|�d�~�f�W�������9��h\�G���u�h�}�8��e����J����\��Y
�����
�
� �g�g��E��Y����^��1��*��a�%�u�h��.����&���� ^����U���6�;�!�9�f�l�L���YӒ��lQ��Q��CҊ�a�i�u�8��l����O����W��S�����|�_�u�u�:��D���&����l��S��D���=�;�}�<�9�9��������l��h]�M���u�<�;�1�6�����&����lV������w�_�u�u�:��C���&����l��S�����:�<�
�0�#�/�����ι�@��R
�����&�2�
�
�"�o�C߁�K����O��N�����b�
� �g�a��E��Yۈ��@��U��G���
�f�c�%�w�2�W�������l
��h_����u�8�
�c�1��D���	���N��P �����
�g�m�%�w�2�W�������l
��h_����u�8�
�b�1��B���	���D�������<�;�1�%��1�(�������
U��G��U���;�1�4�
�8�.�(���M�����RN��W�ߊu�u�8�
�o�;�(��O����[��������!��2�)����&����_9��Q��@���%�u�u�:�;�%�2ߑ�����R��h!��0���9�d�3�
�b�e����_ӄ��_9��r^�����0�!�'���,����&����S��G\����u�8�
�l�1��B���	���D�������8�
�m�3��h�A���Y�ƭ�l��D��ي�|�0�&�u�g�f�W�������l ��\�*��i�u�d�u�?�3�_�������U��
N��*���&�
�#�g�f�t����Y���9F���*���3�
�`�g�'�}�J���[ӑ��]F��Z��M���
�`�c�%�w�}��������EU��N�����e�n�u�u�#�-�Oށ�����9��R��W���"�0�u�!�'�j�(���K����CR������!�9�f�b�w�1����[���F��G1�*���d�a�
�f�k�}��������W��F�U���;�:�d�|�]�}�W���Y����U��B1�Dڊ�d�i�u�!��2����������^�����0�}�
�4�e�e����N�ԓ� O�G����u�u�u�!�'�e�(���K����CW�
N�����2�6�#�6�8�u����ە��]��G1��؊�
� �g�a��n�[��P��ƹF�N�����`�3�
�m�c�-�W��
����\��h�����'�&�/�}�>�3�Ǯ�/����9��h��G��
�f�y�c�~�W�W���Y����^��1��*��m�%�u�h�$�9��������G	��E�����<�;�1�%��1�(�������T��G�C���_�u�u�u�w�)���&����R��G_��Hʦ�1�9�2�6�!�>����������Y�����<�
�<�|�b�t�L�ԜY�Ƹ�C9��Q��Eڊ�d�i�u�'�0�����@Ź��P��N����!�u�|�_�w�}����I���� V��h�I���!�
�:�<��8��������VN��D�����7�4�&�2�����JĹ��J��G�U���!�%�l�
�"�n�Bց�K�����D�����f�3�
�e�f�-�W���Y����\��h��*���_�u�u�8��o����I�Г�F�F����d�'�2�a�f�}����	����@��A_��\�ߊu�u�8�
�d�;�(��I����[�D�����d�'�2�a�o�}����	����@��A_��\�ߊu�u�8�
�c�;�(��H����[��C
�����
�0�!�'�%�.��������V��U1�����
�
� �f�n��E��K����F�C��Lߊ� �f�d�
�e�a�Wǰ�����Q��1��*��e�%�u�:�w�-��������lW�=N��U���
�c�3�
�e�o����D�θ�C9��1����c�u�:�u�'�>�����ד�]ǻN�����b�3�
�g�n�-�W��Q����Q��1����f�u�:�u�'�>�����ד�]ǻN�����m�3�
�f�c�-�W������W��R��D���3�
�f�l�'�u�FϺ�����O��N�����l�
� �f�n��E��Y���D��F��*����&�
�!�"�)����M˹��T9�� [��U���6�;�!�9�d�h�W�������l�N�����3�
�g�g�'�}�J���[ӑ��]F��Y�����&�
�8�
�"�l�F݁�J���F��P ��]���6�;�!�9�f��A�������V�=N��U���
� �d�b��n�K�������]��[��D��!�%�d�
�2��O��B�����h�� ��f�
�g�i�w�l�W����ι�@��R
�����!�3�
�g�e�-�^������]��V�����
�#�g�d�~�}����[����F�B,�����&�
�!� �#�/�(��&����l ��[�*��i�u�!�
�8�4�(�������V��RF�����0�}��6��<��������A��V�����e�`�y�|�l�}�Wϫ�&����R��d�����0�d�m�3��e�E���Y���F�N�����!�%�`�3��j�B���Y����N��h�����
�c�f�%��t�J���^�Ʃ�@�N��U���&�9�!�%�c�;�(��N����9F���*���g�f�
�g�k�}�F������F��P ��]���
��-� ��?��������F�� 1�����a�l�%�|�k�(�����Ϊ�C9��d�����&�9�!�
�6�(�(���H����S��h�\ʰ�&�u�e�n�w�}��������lW��B1�E݊�g�i�u�&�0������ד�F9��W��Fʴ�1�7�8�'�2�o�(�������W��G�U��� �1�'�9� �o����M�Г�F�F����
�0�:�2�9�;�(��I����K	��D�����3�
�g�m�'�t�}���Y����A ��@1�����3�
�a�m�'�}�J�������U��Z�����'�%�f�
��(�E��&���9F������:�
�
� �d�n�(��E����Z��^��*���
�e�a�4�3�)�������� U��G�U��� �1�'�9� �n��������P��N�U¡�%�`�3�
�f�m����Ӗ��9��h��F��
�g�n�u�w�(��������l ��]�*��i�u�&�2�5�)�E�������F��SN�����3�
�f�g�'�t�}���Y����A ��@1�����3�
�f�`�'�}�J�������U��\�����'�%�f�
�e�;�(��H����l�N�����9�"�3�
�f�k����D�ο�T��D�����
�d�e�%�w�3�W�������W��h��G��
�g�n�0�3�?����s