-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�_�&�w�8��������Z��X����_�0�!�!�w��N��Aŀ��l ��O��G���c�
�u�&�w�}�������9F�N��U���u�u�u�u�m�4�������]ǻN��U��� �
���w�g�������F��=N��U���u�<�e����MϷ�����\�\�U���u�u�1� ���#���Y����T��S��A���u�|�_�u�w�2����Y���F��^ �Oʼ�u�&�1�9�0�>�����Ψ�]V��~*��X���:�;�:�e�l�}�W���Yӂ��GF��X�����9�2�6�#�4�2�_�������g.�
�����e�_�u�u�l�8�ϻ�����9l��T�����'�u�'�=�8�}�2��H����lV��G��*���&�c�
�u�$�}�W��T���K�C�X���x�u�:�%�9�3�W��T���K�C�X���x�u�u�6�:�2��������R��Q1�����%�-�
�
�8�9���Y��ƹF�N�����}�u�u�u�w�}�Wϭ�����R9��V��U���u�o�<�u�$�9�������F�N��Uʦ�4�<�
�
�3�)�W���Y����Z�D�����6�#�6�:��l��������l�N��U���u�8�4�<��8��������WF��X�����9�2�6�_�w�}�W���Y�ơ�R��h�� ���!�4�4�u�w�(�W���&����P9��T��]��1�"�!�u�~�}�W���Y����F�R �����:�0�!�_�w�}�Z��T���K�C�X����6�9�&�0�<�W��T���K�C�X�ߊu�u�<�;�;�<��������@��[���ߊu�u�<�;�;�<��������@��[�����6�:�}�d�3�*����P���F��P ��U���#�9�1�o�$�9�������F��P ��U���1�!�u�o�$�9��������G	��]�����:�e�n�7�0�3�W���T���K�C�X���x�x�u�;�#�3�������K�C�X���x�x�u�u�:��B��O����R��G��*ڊ�:�1�%�f��}�W���	����GF��qW�A���
�
�%�3�2�)�G���&���� TǻN�����8�%�}�u�w�}�Wϭ�����R9��V��U���u�h�u�
�!�1��ԜY���F��V��*���1�!�u�u�w�}�IϿ�����l�N��Uʸ�4�<�
�0�"�)���������A���ߊu�u�u�u��%����
����G��VN��Kʧ�!�4�4�u�w�t�}���Y���K�C�X���x�x�x�u�$�4�������K�C�X���x�x�x�u�w�<�������A��d��Uʴ�!�4�4�u�j�u����.����W��X����h�u�e�|� �8�W������N��^ ��"����d�1�"�#�}�W���^���F��F�����u�u�<�e� ��?������\F��
P�� ���|�0�&�u�>�m�}���Y����F�R�����4�4�_�0�3�<��������V]�