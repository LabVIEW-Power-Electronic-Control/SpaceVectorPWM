-- � 2012 National Instruments Corporation.
encrypted

�����'�u���]�.�W���<ݕ��l
��^��D��4�9�_�&�w��2�������l����N���;�<�,�8�g�j�B���&ù��_9��[1����m�
�`�d���O�����A�=N��U��<�u�!�
�8�4�(������F�N�����u�|�_�u�w�g��������T��A�����m�x�d�1� �)�W���s���C\��B�����:�<�
�0�#�/�D���Y�ƨ�D��^��N���;�u�;�<�.�W��������F��U��ʺ�u��l�g��;�G�������lW��D1���
�
��a��}����Yӕ��]��V1�����;�<�;�1�f�}�W�������V�=N��U���;�9�7�6�#�}��������F��S�����|�_�u�u�>�3�Ϯ�����@��R
��@���d�1�"�!�w�t�}����ƓF�V1����u�;�<�;�3�<�L���Yӄ��E�
N�����}�|�_�u�w�����Dӕ��]������� �&�2�0�w�.����Y����@��h��\���&�2�0�u�5�>����Y���l�N��I���!�
�:�<��8����	����]ǑR �����<�0�!�'�l�W�����ƅ�v#��B��<���{�!�
�:�>��F������9��^����b�`�e�
��(�(���&�Ѣ�lW��h]��Dʼ�_�u�u�0�2�4�W�ԜY���F��T��;����n�u�u�w�}�9���*����\��y:��0��u�u�u�u�3�3�(���-����z(��p+�����u�u�u�<�f�
�3���Cӯ��v!��d��U���u�1� �
��	�W���7����aO��N�����u�_�u�u�w�}���Cӯ��`2��{!��6�����}�<�g�
�3���T����|1��xN�N���u�u�u�1�9�}�W���*����|!��h8��!���1�;�
���}�W���6����V�=N��U���u�:�!�o��	�$���5����l0��c!�����
���u�w�}�8���6���l��SN�����n�_�'�=�#�>��������\ ��v^�Gߓ�3�e�8�9�:�1�Fذ�&�޿� S����U���6�8�:�0�#�0�G��L�֪�9��[1����;�
�m�
�b�l�3���A����@l�N��Uʥ�'�u�_�u�w�}�W���Y����z(��c*��:���
����]�}�W���Y���QF��~ ��!�����
����}���Y���F�GN�:���������4���P���F��SN�����0�!�_�_�5�:����YӋ��
Q��q^��E���9�8�9�d�9��O���L�ד�`6��h^��U���6�8�:�0�#�0�G��L�֪�9��[1����;�
�m�
�b�l�3���A��ƹF��X�����}�u�u�u�w�<�J�������F�N����u�<�d�_�w�}�W���Y����\��d�����'�=�!�6�"�8�}��