-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�_�&�w�8��������Z��X����_�0�!�!�w�k�5��:����l ��G1����g�&�d�d�>�W�W�������PF�N��U����u�u�u�w�}�W�������	[�d��U���u������W�������AF��_�U���u�u�1�;���#���Y����T��S��G�ߊu�u�u�u�>�l� ���1����]��R��H��n�u�u�u�w�9����0����	F��C����u�_�u�u�l�}�WϮ����F�N�����u�u�u�;�w�)�(�������P��
��E�����d�1� �)�W���s���F�S��U���u�;�u�!��2����������1��1���d�1�"�!�w�t�}���Y���\��S��U���u�!�
�:�>���������\��XN�N���u�u�u�1�"�}�W����ƿ�W9��P�����:�}�:�!� ��?������\F��=N��U��0�1�0�!�#�f�}�������G����ʺ�u�c��d��;�G�������]�� ��D��<�_�u�u�z�p�Z��T���K�C�6���:�0�!�x�z�p�Z��T���K�CךU���:�%�;�;�w�k�5��:����l��Q��*ڊ�:�1�%�f�w�.�W���Y����\��d��U���u�u�u�&�6�4�(�������F�N��U���;�u�!�
�8�4�L���Y���F������4�!�4�4�w�}�W���Y�ƥ�F��S1�����#�6�:�}�f�9� ���Y����F�N��U���&�4�<�
��+����Y���F���U���
�:�<�n�w�}�W���Y����l��D1�����4�u�u�u�w�}�W���Y����_	��T1�����}�d�1�"�#�}�^�ԜY���F�N�����
�%�'�!�8���������]F��C
�����n�u�u�u�w�}�Wϭ�����\��V�����4�4�u�u�9�}��������E��X��U���;�:�e�n�w�}�W���Y����l��D1�����
�#�9�1�w�}�W���Y����_	��TUךU���u�u�u�u��%����
����G��VN��U��:�!�&�1�;�:��������F��@ ��U���u�u�u�u�~�W�W����Ư�^��R �����u�x�x�x�z�p�Z��T���F��Y�����x�x�x�x�z�p�Z��T���9F�C�4�����:�6�3�W�W�������]��g1��$��&�1�9�2�4�+����Q�ƨ�D��^��O���e�e�d�n�w�}��������r6��p:��U���
�:�<�
�2�)�������\F��T��W��d�w�_�u�w�2����ӧ��|!��N�����2�6�#�6�8�u�W������F��L�E��n�u�u�6�9�)����)����\��C
�����
�0�!�'�c�9� ���Y���F�_�W�ߊu�u�:�&�6�)�6���5����@��[�����6�:�}�u�8�3���Y���V��L�U���6�;�!�;�w��8���Cӕ��l
��^�����'�a�1�"�#�}�^��Y����V�=N��U���&�4�!����W�������T��A�����u�:�;�:�g�}�J���H����l�N�U���c�:�6�1�]�}�W���
����)��r?��Oʦ�1�9�2�6�!�>����Y����G	�N�U��e�e�e�w�]�}�W���
����)��p:��Oʦ�1�9�2�6�!�>����Y����G	�N�U��d�e�e�w�]�}�W���
����)��p+��Oʦ�1�9�2�6�!�>����Y����G	�N�U��d�e�e�w�]�}�W���
����)��{:��Oʦ�1�9�2�6�!�>����Y����G	�N�U��e�d�e�w�]�}�W���
����)��{+��Oʦ�1�9�2�6�!�>����Y����G	�N�U��e�d�e�w�]�}�W���
����)��y+��Oʦ�1�9�2�6�!�>����Y����G	�N�U��d�d�e�w�]�}�W���
����)��b!��Oʦ�1�9�2�6�!�>����Y����G	�N�U��e�e�e�w�]�}�W��T���K�C�X���x��6�9�$�:����T���K�C�X���_�u�u�<�9�1��������\��C
�����n�u�u�&�0�<�W�������F��D�����6�#�6�:��l��������l�N�����u�
�#�9�3�}�W���&����P]ǻN�����9�7�!�4�6�}�Mϭ�����Z��R����u�:�;�:�g�f�W���
����_F��h�����o�&�1�9�0�>�}���Y����R
��G1�����u�u�!�
�8�4�(��������Y��E��u�u�&�2�6�}�(������	F��S1�����_�u�u�<�9�1�������\��C
�����
�0�!�'�`�9� ���Y����Q��Yd��U���x�x�x�x�z�p�Z��T����]��Y�����u�x�x�x�z�p�Z��T���F��r,��D���
�
�%�3�:��(�������9��N�����0�!�8���l�1���&����P��1��*���
�g�u�u�'�/�W���Y���F�N�����
�
�#�9�3�}�W���Y���R9��V��Y���u�u�u�&�6�4�(�������F�N��U��4�!�4�4�]�}�W���Y����Z��h�����u�u�u�u�j�}�(�������F�N�����<�
�
�1�#�}�W���Y���F��C
���ߊu�u�u�u��%��������\��A����u�%�!�4�>�q�W���Y����l��D1�����<�;�!�4�6�}�Iϱ�&����RJǻN��U���
�-�&�'�$�1�(������F������1�_�u�u�w�}�(���
����F
��C
�����u�h�u�
�3�)�}���Y��ƓF�C�X���x�x�x�x�z�p�Zϟ�
����V��C�X���x�x�x�x�z�p�}���Y����R
��N�U��n�u�u�4�#�<����E����Z��`'��=��1�"�!�u�w�c�P���Y����N��^ �H���1�;�
���p�W������[�6��\���'�}�<�e�j�u����&����{K��S�����u�k�r�r�~�}��������9F������1�u�h�r�p�W�W���&����RF�S�����
���x�w�2����I���V������1�;�u�u�w�4�F���=�����Y��E��u��|�u�8�}����Y���W��h9��!���u�:�;�:�g�`�Wȋ�P����_��S��N���u�:�
�#�;�9�K���H��ƹF��X��U���u�h�'�!�6�<�GϺ�����O��=N��U���x�x�x�x�z�p�Z��T�ƃ�P	��C�X���x�x�x�x�z�p�Z��T�����T��Uº�6�1�|�7�0�3�W���Y����R�������u�&�u�u�w�}�W�������r6��r?��Kʺ�
�1�!�u�j��(���s���F�N�����u����j�}�������F��h)�����u�u�u�u�w�5�ϟ�&����X��G1�����i�u���l�}�W���Y�����YN��*���u�k�:�
�3�)�W��6����l�N��U���u�"�0�u���2��Y����W��R��:����_�u�u�w�}�W�������c9��rN��U���!�4�4�i�w��9��Y���F�N������
��u�i�2�(������)��b!�U���u�u�u�u� �8�W������F��h�����h��
��]�}�W���Y����P��d��Uʰ�1�%�:�0�$�W��������G��B��