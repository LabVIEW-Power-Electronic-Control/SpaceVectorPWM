-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�c��m����(���
����GF�N�����9�u�u����;���:���F��h��U���������}���Y����G��T��;ʆ�����]�}�W�������	F��cN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�%�<���6����g"��x)��N���u�<�
�0��1����Y�ƅ�5��h"��<������}�f�9� ���Y����F�^ �����4�
�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���)����W9��N��U���
���
��	�%���Hӂ��]��G�U���<�
�0�
�2�<�G��0�Ɵ�w9��p'��#����u�f�u�8�3���B�����E�����u�u� �u���8���&����|4�_�����:�e�n�u�w�<�(�������\��b:��!�����
����_������\F��d��Uʴ�
�0� �;�e�g�8���*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƭ�l��B��F��������4���:����U��S�����|�_�u�u�'�/����&����|3��d:��9�������w�n�W������]ǻN�����!�'�
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W�������\��yN��1�����|�_�9�f�}������P��RN�����:�u�g��a�i��������@FǻN�����4�!�4�
�8�.�(�������	F��s1��2���o�u�d�n�w�}��������R��X ��*���<�
�u�u���8���Y���A��N�����!�;�u�%���ށ�
����	F��s1��2������u�f�}�������	[�^�E��e�e�e�d�l�}�WϽ�����GF��h=�����3�8�d�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��UךU���:�&�4�!�6��#���J����lT�=��*����
����u�CϺ�����O�
N��E��e�e�e�e�g��}���Y����G����&���!�
�&�
�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��^�N���u�6�;�!�9�}����&����U��N�&���������W��Y����G	�N�U��e�e�e�e�f�m�G��Y����\��V ������&�c�3�:�h�Mύ�=����z%��r-��'���a�1�"�!�w�t�M���I����V��^�E���_�u�u�:�$�<�Ͽ�&����GQ��D��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��[���F��Y�����%��
�!��.�(���Y����)��t1��6���u�d�u�:�9�2�G���D����V��_�E��e�n�u�u�4�3����Y����g9��1����o������!���6���F��@ ��U���o�u�e�e�g�l�G��I���9F������!�4�
��$�l�(���&����`2��{!��6�����u�d�w�2����I����D��^�E��e�e�e�n�w�}��������R��c1��Dۊ�&�
�e�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��UךU���:�&�4�!�6��#���H����^9��T��!�����
����_������\F��T��W��d�e�e�e�g�m�U�ԜY�Ư�]��Y�����
�!�f�3�:�l�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��n�u�u�6�9�)����	����@��h��*��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I���9F������!�4�
��$�l�(���&���5��h"��<������}�c�9� ���Y���F�^�E��e�e�e�w�]�}�W���
������T�����f�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�e�u�W�W�������]��G1�����9�d�d�o���;���:����g)��^�����:�e�u�h�u��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�l�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�F���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�F��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��H����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������wF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����W��L�U���6�;�!�;�w�-��������9��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��_�N���u�6�;�!�9�}��������EW��T��!�����
����_�������V�S��E��u�u�6�;�#�3�W�������l
��h^��U���
���
��	�%���Y����G	�N�U��w�_�u�u�8�.��������]��[�*ٓ�o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��d�d�n�u�w�>�����ƭ�l��D�����f�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��d�e�e�w�]�}�W���
������T�����f�
��o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�d�d�g�f�W�������R��V�����
�#�g��f�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��L�U���6�;�!�;�w�-�������� 9��N��1��������}�A�������V�S��E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-��������9��N�&���������W��Y����G	�N�U��e�e�d�e�f��}���Y����G�������!�9�d�
�a�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��L�U���6�;�!�;�w�-��������9��N�&���������W��Y����G	�N�U��d�d�d�d�g��}���Y����G�������!�9�d�
�b�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��L�U���6�;�!�;�w�-��������lW�=��*����
����u�W������F��L�E��w�_�u�u�8�.��������]��[��F���u��
����2���+����W	��C��\��u�d�e�d�u�W�W�������]��G1�����9�d�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V�=N��U���&�4�!�4��2�����ԓ�\��c*��:���
�����l��������\�^�E��e�e�d�n�w�}��������R��X ��*���g�d�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�d�l�}�WϽ�����GF��h�����#�d�e�o���;���:����g)��_����!�u�|�o�w�m�G��I����]ǻN�����4�!�4�
�8�.�(���M���5��h"��<������}�d�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�d��m�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�N���u�6�;�!�9�}��������EW��q(�Oʆ�������8���H�ƨ�D��^��O���d�d�d�d�g�m�U�ԜY�Ư�]��Y�����;�!�9�d��k�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����W��_�N���u�6�;�!�9�}��������EW��\��U���
���
��	�%���Hӂ��]��G��H���e�e�e�d�g�m�L���YӅ��@��CN��*���&�
�#�g���Mύ�=����z%��r-��'���d�1�"�!�w�t�M���H����W��_�N���u�6�;�!�9�}��������EW��_��U���
���
��	�%���Hӂ��]��G��H���e�e�e�d�g�l�L���YӅ��@��CN��*���&�
�#�g���Mύ�=����z%��r-��'���d�1�"�!�w�t�M���H����W��_�N���u�6�;�!�9�}��������ES��(��3������u�w�	�(���0����p2��F�U���;�:�e�u�j��F��H����W��_�D��d�d�d�d�f�l�F��H����W��_�D��n�u�u�6�9�)����	����@��A_��E��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����A���5��h"��<������}�w�2����I����D��^�E���_�u�u�:�$�<�Ͽ�&����G9��\��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�F��Y����\��V �����:�&�
�#�e��6��*����|!��h8��!���}�d�1�"�#�}�^��Y����W��_�E��u�u�6�;�#�3�W�������l
��1�U����
�����#���Q����\��XN�U��w�e�e�e�f�m�G��Y����\��V �����:�&�
�#�c��1���Y�Ɵ�w9��p'��#����u�g�u�8�3���Y���W��_�D��d�d�d�d�f�l�U�ԜY�Ư�]��Y�����;�!�9�g��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�w�]�}�W���
������T�����d�
��u�w�	�(���0����p2��F�U���;�:�e�u�j��F��H����W�=N��U���&�4�!�4��2�����ԓ�F��d:��9�������w�l�W������F��L�E��e�e�d�w�]�}�W���
������T�����f�
�b�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�d�d�f�f�W�������R��V�����
�#�m�f���Mύ�=����z%��r-��'���b�1�"�!�w�t�M���H����W��_�D��d�n�u�u�4�3����Y����\��h��G��u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��Y����
����m��3���>����v%��eN��Fʱ�"�!�u�|�m�}�G��H����W��_�D��d�d�n�u�w�>�����ƭ�l��D�����m�e�e�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��DҊ���u�u���8���&����|4�Y�����:�e�u�h�u�l�F��H����W��_�����u�:�&�4�#�<�(���
����^��^�U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I���9F������!�4�
�:�$�����@����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
���� T��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��u�u�6�;�#�3�W�������l
��1�U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[��E��������4���Y����\��XN�U��w�e�e�e�g��}���Y����G�������!�9�f�`�m��3���>����v%��eN��U���;�:�e�u�j��G���s���P	��C��U���6�;�!�9�d�k�Mύ�=����z%��r-��'���u�:�;�:�g�}�J���H����F�T�����u�%�6�;�#�1�D��Cӵ��l*��~-��0����}�u�:�9�2�G���D����D��N�����!�;�u�%�4�3����Kƹ��	F��s1��2������u�e�}�������	[�^�E��e�e�e�e�g�m�G��I��ƹF��X �����4�
�:�&��+�(���Y����)��t1��6���u�g�1�"�#�}�^��Y����]ǻN�����4�!�4�
�8�.�(���&����`2��{!��6�����u�g�3�*����P���W��UךU���:�&�4�!�6�����&����F��d:��9�������w�o��������\�^�W�ߊu�u�:�&�6�)��������_��N�&���������W������\F��T��W��w�_�u�u�8�.��������]��[�*��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D�����d�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�d�w�]�}�W���
������T�����f�
�`�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�d�d�f�f�W�������R��V�����
�#�g�d�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�f��k�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�l�F��B�����D��ʴ�
�:�&�
�!�o�D���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�F��H����F�T�����u�%�6�;�#�1�D݁�?����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��H����]ǻN�����4�!�4�
�8�.�(���H���5��h"��<������}�g�9� ���Y���F�^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�g�d�g�$���5����l0��c!��]���:�;�:�e�w�`�U��B�����D��ʴ�
�:�&�
�!��W���-����t/��a+��:���g�1�"�!�w�t�M���I���9F������!�4�
�:�$�����N����u ��N��1��������}�D�������V�S��E��d�d�d�d�f�l�F��H����W��_�N���u�6�;�!�9�}��������EU��^�E��u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��Y�����d�o�����4���:����W��X����u�h�w�d�l�}�WϽ�����GF��h�����#�d�e�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�f��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�l�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s�����Y������3�8�o���;���:����g)��_����!�u�|�o�w�m�G��I����V��UךU���!�'�7�!�w�.�(�������\��C���ߊu�u�!�'�5�)�W���&����W��������3�8�o�$�:����
�Ģ�]�=N��U���;�9�4�
�>�����*����9��Z1�Oʆ�����]�}�W�������C9��P1����u�u����f�W���
����_F��G1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������z0��B��Gۊ�0�
�b�b�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������C9��P1������&�b�3�:�k�Mύ�=����z%��N�����4�u�%�&�0�?���Y�Ǝ�|*��yUךU���<�;�9�2�'�;�(��&���5��h"��<������}�f�9� ���Y����F�D������-��,�"��Fׁ�����T�=��*����
����u�FϺ�����O��N�����4�u�&�0��8�(��N����g"��x)��*�����}�u�8�3���B�����Y�����<�
�&�$���ׁ�
����	F��s1��2���_�u�u�<�9�1��������W9��T��:����n�u�u�$�:��������l ��Y�����u��
����2���+������Y��E��u�u�&�2�6�}����J����lU�� N�&���������W��Y����G	�UךU���<�;�9�!�'�k����N˹��\��c*��:���
�����}�������9F������!�%�c�'�0�n�@���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��(�����m�
�g�o���;���:����g)��_����!�u�|�_�w�}����Ӡ��A��Y�U����
�����#���Q����\��XN�N���u�&�2�4�w��9���:���� _��G\��U���
���
��	�%���Y����G	�UךU���<�;�9����9�������
T�=��*����
����u�W������]ǻN�����9�!�%�a��(�C���	����`2��{!��6�����u�`�3�*����P���F��P ��U���
�f�'�2�d�d�W���-����t/��a+��:���`�1�"�!�w�t�}���Y����R
��T�����`�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����l��h]�F��������4���Y����\��XN�N���u�&�2�4�w�.����&����R��N�&���������W������\F��d��Uʦ�2�4�u�&�2��(���&����\��c*��:���
�����}�������9F������!�%�f�
�"�h�E���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����m�'�2�f�f�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������hZ�����b�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����T��R	��M���o������!���6�����Y��E��u�u�&�2�6�}����HĹ��lS��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�#�-�F�������U��N��1��������}�F�������V�=N��U���;�9�!�%�f�e����Hù��\��c*��:���
�����j��������l�N�����u�8�
�d��8�(��L����g"��x)��*�����}�b�3�*����P���F��P ��U���d�3�
�f��n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h_�����m�e�o����0���/����aF�
�����e�n�u�u�$�:����&¹��lQ��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u������A���5��h"��<������}�w�2����I��ƹF��^	��ʦ�9�!�%�l�1��Fف�J����g"��x)��*�����}�b�3�*����P���F��P ��U���
�8�g�
�2��O��Cӵ��l*��~-��0����}�b�1� �)�W���s���@��V�����8�f�
� �`�m����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���f�
�0�
�o�h�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�`�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��B���2�f�c�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӏ��CT��B1�G���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����K����lU��N�&���������W������\F��d��Uʦ�2�4�u�8��m����I˹��\��c*��:���
�����}�������9F������!�%�c�
�2��O��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
�9�
�;�$�l�ށ�����l��N��1��������}�GϺ�����O��N�����4�u�4�2�e�<��������ZW��R	��M��o������!���6�����Y��E��u�u�&�2�6�}����H����l	��D1��ۊ� �l�a�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������R��1�����0�
�
�d�%�:�D��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����d�4�9�/�%�.�E���&����V��G]��U���
���
��	�%���Y����G	�UךU���<�;�9��9�8�(���&����@9��^_�����m�f�o����0���/����aF�
�����e�n�u�u�$�:����&�Г�9��h_�C���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1���&�ד�V��W�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��<�E�������S��N�&���������W��Y����G	�UךU���<�;�9�%��1�(ہ�����U�=��*����
����u�DϺ�����O��N�����4�u�%�&�0�>����-����l ��hV��U���
���n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��@�����
�0�
�l�g�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��\�� ��`�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����T��R	��L��o������!���6�����Y��E��u�u�&�2�6�}��������A	��Q��@���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϻ�����l��X�����l�a�o����0���/����aF�
�����e�n�u�u�$�:��������W9��R�� ��d�
�f�o���;���:����g)��^�����:�e�n�u�w�.����Y����G��X ��*���
�l�l�o���;���:����g)��^�����:�e�n�u�w�.����Y����VW��[�����g�<�d�
�"�l�E܁�K����g"��x)��*�����}�u�8�3���B�����Y��'���0�
�9�
�9�.�E���Hǹ��T9��Z��U���
���
��	�%���Y����G	�UךU���<�;�9�%��1�(�������U��N�&���������W��Y����G	�UךU���<�;�9�%��1�(�������
U��N��1��������}�F�������V�=N��U���;�9�:�0�1�2�(ށ�����9��T��!�����
����_�������V�=N��U���;�9�:�0�1�2�(ށ�����P�=��*����
����u�W������]ǻN�����9� �1�'�;�*�F���&����l��N��1��������}�GϺ�����O��N�����4�u�;�0�1�2�(ށ�����W�=��*����
����u�W������]ǻN�����9�7�8�'�2����@����\��c*��:���
�����}�������9F������7�8�'�0��8�(��N����g"��x)��*�����}�u�8�3���B�����Y�����9�
�c�3��m�A���Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����9�
�c�'�0�n�A���Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N��*���
�&�$���)�G������5��h"��<��u�u�&�2�6�}��������lW��T��:����n�u�u�$�:��������9��P1�B���u��
����2���+����W	��C��\�ߊu�u�<�;�;�.��������W��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�>�3��������P�=��*����
����u�W������]ǻN�����9�%��9��m����K�Փ�F��d:��9�������w�o�W������]ǻN�����9�%��9��m����J����	F��s1��2������u�e�}�������9F������;�"�<�;�>��(���K����CU�=��*����
����u�W������]ǻN�����9�;�"�<�9�4�(݁�����
V�=��*����
����u�W������]ǻN�����9�6�'�,�1��E���	����`2��{!��6�����u�e�3�*����P���F��P ��U���'�
�0�
�n�j�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[�����'�&�g�3��o�F���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����0�
�0�:������I���5��h"��<������}�w�2����I��ƹF��^	��ʥ��9�
�d�1��D���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʥ��9�
�d�%�:�C��Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����<�
�&�$����������F��d:��9����_�u�u�>�3�Ͽ�&����Q��V�Oʗ����_�w�}����ӏ��CU��B1�G؊�g�o�����4���:����V��X����n�u�u�&�0�<�W���	����T9��]��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�e�(���K����CT�=��*����
����u�W������]ǻN�����9�!�%�m��8�(��A����g"��x)��*�����}�u�8�3���B�����Y�����m�
� �g�c��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��M؊�0�
�e�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G[�����a�m�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��^�����e�e�o����0���/����aF�
�����e�n�u�u�$�:��������CS��Q��A���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����T��R	��E��o������!���6�����Y��E��u�u�&�2�6�}��������U��W�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	�Փ�V��Z�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�'�.��������l��1����u�u��
���L���Yӕ��]��V�����1�
�e�u�w��;���B�����Y�����!�%�a�3��h�B���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�`�
�0��m�A��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��B,�����&�
�!� �#�/�(��&����P��G]��U���
���
��	�%���Y����G	�UךU���<�;�9� ��.�4���&����P��R1�M���2�a�c�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��]��h_�����e�d�o����0���/����aF�
�����e�n�u�u�$�:����&����lS��E��A��u�u��
���(���-��� W��X����n�u�u�&�0�<�W����ד�V��V�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��C؁�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��i�(���&����\��c*��:���
�����m��������l�N�����u�8�
�a��8�(��K����g"��x)��*�����}�u�8�3���B�����Y�����d�l�'�2�c�d�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��@ۊ�0�
�d�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƽ�a��[��*���'�2�a�e�w�}�#���6����e#��x<��Dʱ�"�!�u�|�]�}�W�������l4��B��D���2�a�d�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��]��h\�����d�m�o����0���/����aF�
�����e�n�u�u�$�:����&����lS��E��A��u�u��
���(���-��� W��X����n�u�u�&�0�<�W����ԓ�V��\�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��Bہ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��h�(���&����\��c*��:���
�����m��������l�N�����u�8�
�`��8�(��@����g"��x)��*�����}�u�8�3���B�����Y�����d�c�'�2�c�i�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��@Ҋ�0�
�d�l�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƽ�a��[��*���
�d�a�o���;���:����g)��_�����:�e�n�u�w�.����Y����@��hZ�����d�l�o����0���/����aF�
�����e�n�u�u�$�:��������
9��P1�C���u��
����2���+����W	��C��\�ߊu�u�<�;�;�-�!���&����l ��^�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������_��R	��D��o������!���6���F��@ ��U���_�u�u�<�9�1��������V��c1��Dي�&�
�g�o���;���:���F��P ��U���&�2�7�1�e�d�MϜ�6����l�N�����u�
�4�g�b����K˹��\��c*��:���
�����l��������l�N�����u�
�4�g�b�����H���5��h"��<������}�f�9� ���Y����F�D������6�
�4�2���������W��1��*��g�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G9��D�����!�'�
�b��l����M����	F��s1��2������u�d�}�������9F������4�
�<�
�$�,�$����ғ�@��N�&������_�w�}����Ӈ��@��U
��G��o�����W�W���������T������'�6� �2�l�O�������R��N�&���������W��Y����G	�UךU���<�;�9�<��)�4���&����P��R1�M���'�2�a�m�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����Z*��C1�����!� �!�'��e�(ց�����9��T��!�����
����_������\F��d��Uʦ�2�4�u��4�����*����G��h_�*ӊ�0�
�d�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������V��Q��A���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϭ�˹��T9��V��U���
���
��	�%���Y����G	�UךU���<�;�9�<��4�1���5����_��Q��A���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ͽ�&����P��h=����
�&�
�a�m��3���>����F�D�����%�&�2�7�3�o�@��;����r(��N�����4�u�'�
�#���������9��R1��D���
�c�f�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����V��T��*���f�`�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƭ�A9��h(��*���%�g�a�g�2�m�D���&����l��N��1��������}�D�������V�=N��U���;�9�4�'�;���������R��h��*ߊ� �f�a�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��3����:�
�e���(ށ�&����S��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%���������C9��1�����f�3�
�c�f�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��V�����:�
�:�%�e�i�E���H�ӓ�F9��Y��F��������4���Y����W	��C��\�ߊu�u�<�;�;�>�(���<����G��h\�*���
�0�
�a�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����P
��y*��4���0�8�g�a�2�m����K���5��h"��<������}�f�9� ���Y����F�D�����'�
�!��%�����Iǹ��V9��1����a�o�����4���:����U��S�����|�_�u�u�>�3�Ͽ�����u	��{��*��
�
�
�
�2��@���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*������0�:�o�C���H����lT��T��!�����
����_������\F��d��Uʦ�2�4�u�9���/�������U��R1�����g�b�o����0���/����aF�N�����u�|�_�u�w�4��������l ��h"�����'�2�f�m�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƫ�C9��h]�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������9��T��!�����
����_������\F��d��Uʦ�2�4�u�'��(�D���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʲ�%�3�
�g��l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��h�����3�
�f�
�g�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������D�����3�
�f�
�g�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������D�����
�f�
�d�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������A��a1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������^��h��F���%�u�u����>���<����N��
�����e�n�u�u�$�:��������U��Z��D��������4���Y����W	��C��\�ߊu�u�<�;�;�)��������9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��k����@Ź��\��c*��:���
�����l��������l�N�����u�8�
�a�1��Gׁ�H����g"��x)��*�����}�u�8�3���B�����Y�����d�
� �a�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h�����d�
�g�o���;���:����g)��[�����:�e�n�u�w�.����Y����V��V�����
� �a�c�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�����c�
�g�o���;���:����g)��_����!�u�|�_�w�}����Ӓ��lT��Q��Fފ�g�o�����4���:����W��S�����|�_�u�u�>�3�Ϫ�	����U��^��A��������4���Y����W	��C��\�ߊu�u�<�;�;�9��������U��[��D��������4���Y����W	��C��\�ߊu�u�<�;�;�4����&¹��lR��h�Oʆ�������8���O�ƨ�D��^����u�<�;�9�2�-����/�ד�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��l�(���M�ԓ�F��d:��9�������w�h�W������]ǻN�����9�!�%�f��(�C���	����`2��{!��6�����u�`�w�2����I��ƹF��^	��ʥ��&�9�
��(�B���	����`2��{!��6�����u�`�w�2����I��ƹF��^	��ʸ�;��f�3��m�(��Cӵ��l*��~-��0����}�f�1� �)�W���s���@��V�����d�
� �a�g�-�W���-����t/��a+��:���c�u�:�;�8�m�L���Yӕ��]��q\��*���`�m�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ɲ�r(��y-��*���`�a�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lU��Q��Aڊ�g�o�����4���:����W��S�����|�_�u�u�>�3�Ϫ�	����U��X��G��������4���Y����W	��C��\�ߊu�u�<�;�;�.�(���&¹��lS��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�:�3�!�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�=�6�)�F���
����lS��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�#�-�Cځ�����l��N��1��������}�B�������V�=N��U���;�9�!�%�c����I����	F��s1��2������u�b�}�������9F������!�%�d�c�1��@߁�H����g"��x)��*�����}�b�3�*����P���F��P ��U���
�b�3�
�g��F��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���3�
�e�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h[�����g�
�g�o���;���:����g)��_����!�u�|�_�w�}����Ӓ��lP��T��*���c�c�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��C���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����l ��]�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����T��N�&���������W��Y����G	�UךU���<�;�9�!�'�l�G���&����CW�=��*����
����u�W������]ǻN�����9�!�%�`��(�A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���%�
� �c�o�-�W���-����t/��a+��:���`�1�"�!�w�t�}���Y����R
��Z��Gۊ� �c�a�%�w�}�#���6����e#��x<��@ʱ�"�!�u�|�]�}�W�������^��\�� ��g�%�u�u���8���&����|4�]�����:�e�n�u�w�.����Y����T��Q��M܊�g�o�����4���:����S��S�����|�_�u�u�>�3�Ϫ�	����l ��W�����u��
����2���+������Y��E��u�u�&�2�6�}�(�������l ��W�����u��
����2���+������Y��E��u�u�&�2�6�}����J����R��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�h�(���N�ғ�F��d:��9�������w�m��������l�N�����u�8�
�d�1��Aہ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�e�3��o�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����l�3�
�f��i�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��Z�����a�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����R��B1�E���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����HĹ��@��V�����`�
�f�o���;���:����g)��_����!�u�|�_�w�}����Ӄ��l0��h��A���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l �� X�����u��
����2���+������Y��E��u�u�&�2�6�}����Jù��lQ��h�Oʆ�������8���H�ƨ�D��^����u�<�;�9�'�.�(ށ�����l��N��1��������}�F�������V�=N��U���;�9�%�&�����A����	F��s1��2������u�f�}�������9F������!�%�d�g�1��Fہ�J����g"��x)��*�����}�u�8�3���B�����Y�����
�
�4�!�1��Nہ�H����g"��x)��*�����}�d�3�*����P���F��P ��U���
�d�3�
�e��F��*����|!��h8��!���}�f�1�"�#�}�^�ԜY�ƿ�T����*���3�
�f�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W�������
��1��*��
�d�o����0���/����aF�
�����e�n�u�u�$�:�����ԓ�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�(���A�ԓ�F��d:��9�������w�m��������l�N�����u�8�
�f��(�O���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�a�3�
�a��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��E��*���m�g�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӗ��9��T��*���m�a�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��M���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l0��h��M���%�u�u����>���<����N��
�����e�n�u�u�$�:����&����U��^��G��������4���Y����W	��C��\�ߊu�u�<�;�;�2�(����ד�9��hV�*��o������!���6�����Y��E��u�u�&�2�6�}����K����l	��D1�����l�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����VW��[�����f�3�
�a��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���l�g�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӵ��T��V�����&�g�3�
�e��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��e��ۊ�9�
�0�:�����O����	F��s1��2������u�g�9� ���Y����F�D�����8�
�b�;�#�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�c�
� �n�m����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���f�
� �l�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����
� �l�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W�������	��T��Lي�d�3�
�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��Y	��*���
�;�&�g�1��Fف�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�e�3��j�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��Lߊ�d�3�
�`��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��V��D���
�f�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��GZ�����l�
�f�o���;���:����g)��^�����:�e�n�u�w�.����Y����U��Q��E���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����V��h�Oʆ�������8���L�ƨ�D��^����u�<�;�9�'�����&Ź��lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�<�(���&����U��G\��U���
���
��	�%���Jӂ��]��G�U���&�2�4�u�:��(���H����CT�=��*����
����u�FϺ�����O��N�����4�u�8�
��(�F��&���5��h"��<������}�f�9� ���Y����F�D�����=�4�!�3��m�A���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y������3�
�e�n�-�W���-����t/��a+��:���`�u�:�;�8�m�L���Yӕ��]��D�����4�!�3�
�g�n����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����3�
�e�m�'�}�W���&����p9��t:��U���u�:�;�:�g�f�W���
����_F��G1�����e�g�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��h��D��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������9��h_�L���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&�ד�F9��]��G��������4���Y����W	��C��\�ߊu�u�<�;�;�)��������P��N�&���������W������\F��d��Uʦ�2�4�u�8��n����I�ޓ�F��d:��9�������w�o�W������]ǻN�����9�%�g�3��l�E���Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����d�
� �d�d��E��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���6�&�
� �f�i�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����g�3�
�d�f�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��M���
�d�c�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��1��*��c�%�u�u���8���&����|4�]�����:�e�n�u�w�.����Y����W��B1�Cӊ�g�o�����4���:����S��S�����|�_�u�u�>�3�Ϫ�	����U��Y�����u��
����2���+������Y��E��u�u�&�2�6�}�(�������l ��_�*��o������!���6��� F��@ ��U���_�u�u�<�9�1����Hƹ��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Fׁ�����9��T��!�����
����_�������V�=N��U���;�9�%��;��(���H����CU�=��*����
����u�DϺ�����O��N�����4�u�8�
�a�;�(��N����	F��s1��2������u�g�9� ���Y����F�D�����
� �d�l��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��^1�����g�d�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӗ��U��[�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�,�(�������l ��\�*��o������!���6�����Y��E��u�u�&�2�6�}����I����T��h�Oʆ�������8���K�ƨ�D��^����u�<�;�9�'��݁�&����T��G\��U���
���
��	�%���Jӂ��]��G�U���&�2�4�u�:��(���H����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'����Mʹ��\��c*��:���
�����}�������9F������&�9�!�%��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�c�
� �f�d�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�d�3�
�e�m����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���f�3�
�g�f�-�W���-����t/��a+��:���g�u�:�;�8�m�L���Yӕ��]��D�����f�3�
�g�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����
� �d�m��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�g�c�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��[1�����3�
�g�a�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h[�� ��m�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����G�� 1��*��l�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������9��h_�L���u�u��
���(���-���U��X����n�u�u�&�0�<�W���&����9��h_�C���u�u��
���(���-���U��X����n�u�u�&�0�<�W���&�ԓ�F9��]��F��������4���Y����\��XN�N���u�&�2�4�w�0�D�������T��Q��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	¹��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'�.�(���H����CT�=��*����
����u�FϺ�����O��N�����4�u�:�g�1��D���	����`2��{!��6�����u�d�w�2����I��ƹF��^	��ʡ�%�d�c�3��n�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����6�&�
� �f�n�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����a�3�
�f�`�-�W���-����t/��a+��:���`�u�:�;�8�m�L���Yӕ��]��C��G܊� �d�m�
�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W�������
��Q��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϭ�����U��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:�o����J�ד�F��d:��9�������w�m��������l�N�����u�8�
�e��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�g�
� �f�l�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��ۊ� �d�d�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����C	��h�����
�f�`�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����G��W�� ��g�
�d�o���;���:����g)��[����!�u�|�_�w�}����Ӵ��T��a1�����a�f�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƾ�e9��h_�L���u�u��
���(���-���U��X����n�u�u�&�0�<�W�������9��Q��A���%�u�u����>���<����N��S�����|�_�u�u�>�3�ό�����R
��X ��*���d�a�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�d�<�3��i�F���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����d�4�9�:�2��(���H����CT�=��*����
����u�W������]ǻN�����9�!�%�f��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʇ�;�0�
�9��8��������9��T��!�����
����_�������V�=N��U���;�9��;�2���������9��h_�@���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Kʹ��G9��h_�B���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����J¹��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����A����S��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����W��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�:��2��������R��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�6�:�F�������@9��h_�@���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l ��[�*��o������!���6�����Y��E��u�u�&�2�6�}�(�������S��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��e����&����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�o�(���H����CU�=��*����
����u�W������]ǻN�����9�6�'�,�f�4����J�ӓ�F��d:��9�������w�m��������l�N�����u�4�2�d�6�1����&����U��]�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�����&����I��D1�����
�`�l�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���
� �d�c��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G]�� ��b�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����J9��Y�����
�`�b�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������R��1�����0�
�
�:�����A����\��c*��:���
�����}�������9F������!�%�d�g�1��A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���0�2�l�
��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʇ�;�0�
�9��3��������l ��[�*��o������!���6�����Y��E��u�u�&�2�6�}�(�������P��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�����Kʹ��\��c*��:���
�����j��������l�N�����u�
�4�g�n�;�(��O����	F��s1��2������u�f�}�������9F������!�%�d�b�1��A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�d�3�
�a�i����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������2�
�
� �f�h�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
� �d�c��l�Mύ�=����z%��r-��'���b�1�"�!�w�t�}���Y����R
��h8��G���3�
�c�m�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�C���
�c�g�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���d�m�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G]�����c�a�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��[�� ��e�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����G��1��*��b�%�u�u���8���&����|4�Y�����:�e�n�u�w�.����Y����G��1��*��`�%�u�u���8���&����|4�Y�����:�e�n�u�w�.����Y����T��Q��C���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����W��E	��*���d�d�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�CQ��B1�Gފ�g�o�����4���:����V��X����n�u�u�&�0�<�W�������ZW��B1�Fڊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����R��X�� ��`�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����l ��Y�*��o������!���6�����Y��E��u�u�&�2�6�}����&¹��G9��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������l��h�����;�!�<�
�"�l�A؁�K����g"��x)��*�����}�u�8�3���B�����Y�����'�0�l�<��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʇ�;�0�
�9��3��������9��h_�M���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1�%���¹��_9��R��*���d�
� �d�n��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��S�����:�0�
�
�"�l�O܁�J����g"��x)��*�����}�u�8�3���B�����Y�����!�%�g�3��e�F���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����2�7�!�d�1��@���	����`2��{!��6�����u�e�3�*����P���F��P ��U���d�
� �d�f��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����a�3�
�m�d�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��L���
�b�`�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���d�d�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƨ�_��S1�����d�3�
�b�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R�����0�:�
�
�8����Jƹ��\��c*��:���
�����}�������9F������1�9�!�1�-�/��������9��h_�D���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������9��h_�C���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����N¹��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�3�1��������9��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������V_��S�����
�d�3�
�o�n����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������&�2�
�
�"�l�E؁�J����g"��x)��*�����}�u�8�3���B�����Y�����'�0�b�<��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʦ�2�
�&�<�9�l��������W��N�&���������W������\F��d��Uʦ�2�4�u�8�f����AĹ��\��c*��:���
�����}�������9F������&�9�!�%�e�;�(��M����	F��s1��2������u�g�9� ���Y����F�D�����8�a�3�
�n�i����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���g�
� �d�e��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��Fي� �d�l�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��F���
�l�l�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��R
�����
�:�
� �f�n�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����1�/�'�&�g�3��������W��N�&���������W������\F��d��Uʦ�2�4�u�'�2�:�(�������9��T��!�����
����_�������V�=N��U���;�9�!�%�d����L¹��\��c*��:���
�����}�������9F������1�9�!�1�8�8�(߁�&����
V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�7�:�/��������T��^1��*��g�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����R��P �� ��g�
�f�o���;���:����g)��^�����:�e�n�u�w�.����Y����A�� 1�����l�b�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӓ��V��X�� ��b�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����U
��h��D���
�g�o����0���/����aF�
�����e�n�u�u�$�:��������@��Y1�����
�l�`�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��Q��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϼ�����l��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}�(���K�ӓ�F9��^��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.����	�ѓ�V��P�����e�l�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��[�� ��g�
�f�o���;���:����g)��\����!�u�|�_�w�}����ӄ��V��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CT��Q��E���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	Ź��lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����A����V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u��<�E�������F9��]��F��������4���Y����W	��C��\�ߊu�u�<�;�;�.����	�Г�F9��]��F��������4���Y����W	��C��\�ߊu�u�<�;�;�?��������9��h\�A���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Nù��lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'��݁�&����Q��G]��U���
���
��	�%���Nӂ��]��G�U���&�2�4�u�2����J����\��Y1��*��f�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��h��G��
�f�o����0���/����aF� N�����u�|�_�u�w�4����
����^��h��G��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������U��^�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	�ޓ�F9��Z��G��������4���Y����\��XN�N���u�&�2�4�w�����Hù��K9��h\�M���u�u��
���(���-���Q��X����n�u�u�&�0�<�W���&����9��h\�B���u�u��
���(���-���Q��X����n�u�u�&�0�<�W���&����9��1�����d�l�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�e��h\�����d�l�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�e��h\�����d�l�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��1��*��d�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������W��B1�Mӊ�f�o�����4���:����V��X����n�u�u�&�0�<�W���&����Q��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�'�>�4�(���K����CT�=��*����
����u�W������]ǻN�����9�$�<�
�"�o�A܁�J����g"��x)��*�����}�u�8�3���B�����Y�����&�<�;�`�1��E���	����`2��{!��6�����u�e�3�*����P���F��P ��U���4�g�g�
�"�o�B܁�M����g"��x)��*�����}�f�3�*����P���F��P ��U���
�a�3�
�e�d����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N����e�3�
�d�f�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��@���
�g�b�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������l4��B��Dފ�:�
� �g�d��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��Y�����,�3�
�g�b�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��F���
�g�g�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������K��u=�� ���7�:� �0��1���&����lT�� 1��U����
�����#���Q����\��XN�N���u�&�2�4�w�����&����^��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�7�:�/����&����_��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�j�(���K����CT�=��*����
����u�W������]ǻN�����9�%�f�
��(�E��&���5��h"��<������}�w�2����I��ƹF��^	��ʷ�8�'�0�e�3�0����&����lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�E܁�����R��B1�EҊ�g�o�����4���:����V��X����n�u�u�&�0�<�W�������D9��Q��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϱ�����D9��Q��G���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	�Փ�F9��[��G��������4���Y����\��XN�N���u�&�2�4�w�/����&����l ��]�*��o������!���6�����Y��E��u�u�&�2�6�}��������9��C1��*��e�%�u�u���8���&����|4�N�����u�|�_�u�w�4����	����9��h��*���g�f�
�f�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������l0��1�����f�f�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƹ�C9��1��*��m�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������9��h\�G���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����8����F��U�� ����9�0�l�����N˹��\��c*��:���
�����n��������l�N�����u�-�
��/�(�(�������l0��B��B���3�
�g�g�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��&���!��&�9�#�����&�ߓ�l ��]�*��o������!���6��� F��@ ��U���_�u�u�<�9�1��������
T��N�&���������W������\F��d��Uʦ�2�4�u�:�;�%�2�������R��h!��0���9�&�3�
�d�e����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T���������!��2�)����&����_9��Q��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϼ�����vV��C1�����'��
�$�6��(���K����CT�=��*����
����u�W������]ǻN�����9�!�%�d�c�;�(��M����	F��s1��2������u�f�9� ���Y����F�D�����8�
�m�3��i�C���Y�Ɵ�w9��p'��#����u�g�1� �)�W���s���@��V�����3�
�a�m�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��Aӊ� �g�`�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����Z��Y����� �g�b�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G�� W�� ��f�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����G��1��*��c�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��1�����4�
� �g�a��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����m�
�0�:�0�3����M�ޓ�F��d:��9�������w�m��������l�N�����u�-�
�:�2�)����Mù��U��^�����u��
����2���+������Y��E��u�u�&�2�6�}��������V��^��#���
�`�l�%�w�}�#���6����e#��x<��G���:�;�:�e�l�}�Wϭ�����U��Y��*���8�`�d��1��B���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʺ�
�:�1�3��h�N���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����9�3�
�`�c�-�W���-����t/��a+��:���g�u�:�;�8�m�L���Yӕ��]��X�����
� �g�a��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h��؊� �g�`�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����]��R�����`�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�C9��S�����a�b��3��h�D���Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����0�f�3�
�b�j����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N�����`�3�
�`�e�-�W���-����t/��a+��:���g�u�:�;�8�m�L���Yӕ��]��Y�����3�
�`�`�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��@=��L���
�c�c�%�w�}�#���6����e#��x<��G���:�;�:�e�l�}�Wϭ�����]��R�G���&�
� �g�f��F��*����|!��h8��!���}�a�1�"�#�}�^�ԜY�ƿ�T�� ��&���
� �g�g��n�Mύ�=����z%��r-��'���a�1�"�!�w�t�}���Y����R
��R��؊� �g�d�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��@ߊ� �g�f�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����C9��Q��@���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����Q��B1�@ފ�f�o�����4���:����T��X����n�u�u�&�0�<�W���&����9��h\�C���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������U��]�����u��
����2���+������Y��E��u�u�&�2�6�}�(���K�ѓ�F9��V��F��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����Q��G_��U���
���
��	�%���Lӂ��]��G�U���&�2�4�u�:��C���&����l��N��1��������}�E�������V�=N��U���;�9�%��;��(�������
V��N�&���������W��Y����G	�UךU���<�;�9�%��1�(�������_��N�&���������W��Y����G	�UךU���<�;�9�!�'�e�(���K����CW�=��*����
����u�BϺ�����O��N�����4�u�8�
�a�;�(��A����	F��s1��2������u�e�}�������9F������'��a�3��k�O���Y�Ɵ�w9��p'��#����u�g�u�8�3���B�����Y�����-� ���#���������9��Q��B���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l ��Y�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������J)��h#�����,�d�a��1��@���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʧ��`�3�
�a�o����Y����)��t1��6���u�g�u�:�9�2�G��Y����Z��[N����� ���!��1����&����e9��h\�C���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����g��C1�����9�
�g�
��(�E��&���5��h"��<������}�b�9� ���Y����F�D�����-�
���.�(�(�������lW��h8�� ��e�
�g�o���;���:����g)��[����!�u�|�_�w�}����Ӏ��l��{:�� ��� �!�%�,�f�j�!���&����l��N��1��������}�B�������V�=N��U���;�9�'�f�1��O���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�f�3�
�o�n����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������2�
�
� �e�e�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
� �g�l��l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��h8��G���
� �g�l��o�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��R�����!�f�3�
�n�o����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���3�
�l�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������E��*���g�d�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�`�3�
�n�k����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T��<�����4�9�/�'�$�i����@�ד�F��d:��9�������w�m��������l�N�����u�4�2�g�6�1����&����lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�N݁�����9��T��!�����
����_�������V�=N��U���;�9�%�a��l����@�ߓ�F��d:��9�������w�m��������l�N�����u�0�0�0��8����&����
U��G]��U���
���
��	�%���Y����G	�UךU���<�;�9�%�9�)�ށ�����
9��T��!�����
����_�������V�=N��U���;�9�7�8�%�8�܁�����9��T��!�����
����_�������V�=N��U���;�9�!�%�n����A¹��\��c*��:���
�����}�������9F������1�9�!�1�8�8�(݁�����9��T��!�����
����_�������V�=N��U���;�9�%�f��l����@�Փ�F��d:��9�������w�m��������l�N�����u�'�0�2�c���������9��h\�G���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Kƹ��^	��V �� ��l�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����9��h]�A���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������lU��B1�Dڊ�g�o�����4���:����V��X����n�u�u�&�0�<�W�������lU��B1�M܊�g�o�����4���:����V��X����n�u�u�&�0�<�W���Hƹ��lU��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�5�0��������U��_�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�(��������l��h��F��
�g�o����0���/����aF�
�����e�n�u�u�$�:����&����lT��h��*���f�f�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������l0��1��DҊ� �f�a�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��F���
�g�o����0���/����aF�
�����e�n�u�u�$�:����&����l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}����
����
9��h]�B���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����@ǹ��lU��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�����L����lU��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�8��������l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}����L���� V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�6�/�(݁�����9��T��!�����
����_�������V�=N��U���;�9��;�2���������l ��_�*��o������!���6�����Y��E��u�u�&�2�6�}����H����l��X��*���f�d�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�a�3�
�f�m����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���3�
�d�f�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������1��*���f�g�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƨ�_��S1�����a�3�
�d�b�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h ��*���3�
�d�m�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������R��*���3�
�d�a�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������hW�����d�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӂ��V��h�����3�
�d�a�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������1��*���f�a�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ʈ�^��RZ�����'�4�
�g�1��F���	����`2��{!��6�����u�e�3�*����P���F��P ��U���f�b�1�8�%�<�(���J����CT�=��*����
����u�W������]ǻN�����9�!�%�c�1��F���	����`2��{!��6�����u�e�3�*����P���F��P ��U���0�3�:�
��(�D��&���5��h"��<������}�w�2����I��ƹF��^	��ʺ�0�3�:�
��(�D��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�b�3�
�e�m����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������
�
�a�3��l�C���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����3�:�
�
�8����IŹ��\��c*��:���
�����}�������9F������%��9�
�g���������9��T��!�����
����_������\F��d��Uʦ�2�4�u�
�6�o�D��&����T��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�:�l�(���J����CT�=��*����
����u�FϺ�����O��N�����4�u��;�3�����H�֓�F9��^��G��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����R��GZ��U���
���
��	�%���Iӂ��]��G�U���&�2�4�u��>�(�������F��E��BҊ�
� �f�`��l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��{1��*���0��'�6�"�8�F���Hù��lU��1��U����
�����#���Q����\��XN�N���u�&�2�4�w���������G��C��*��
�
� �f�a��E��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���3�
�g�l�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������T������'�6� �2�l�F���&����l��N��1��������}�D�������V�=N��U���;�9�!�%�f�m����K�ғ�F��d:��9�������w�m��������l�N�����u�0�
�8�b����H˹��\��c*��:���
�����}�������9F������&�9�!�%�n�;�(��M����	F��s1��2������u�g�9� ���Y����F�D������6�
�4�2���������W��h��F��
�f�o����0���/����aF�N�����u�|�_�u�w�4����
����^�� 1�����4�
� �f�d��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��D���3�
�g�l�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��Cڊ� �f�a�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��D���
�f�e�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������9��h-�����'�6� �0�f�l�E���&����l��N��1��������}�D�������V�=N��U���;�9�&�9�#�-�@ہ�����R��B1�Cފ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����U��V�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	�ԓ�F9�� ^��G��������4���Y����\��XN�N���u�&�2�4�w�8�(���O����lU��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�>�����
����A��B��D���f�3�
�f�a�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��^"�����&�
�!� �#�/�(��&����_��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u��>�(�������F��E��BҊ�
� �f�l��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��{1��*���0��'�6�"�8�F���K���� U��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�>�����
����A��B��D���f�3�
�a�a�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��^"�����&�
�!� �#�/�(��&����lU��1��U����
�����#���Q����\��XN�N���u�&�2�4�w���������G��C��*��
� �f�g��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��{1��*���0��'�6�"�8�F���M���� R��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�>�����
����A��B��D���`�3�
�a�o�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��D�����3�
�a�d�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��G���
�a�f�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������9��h-�����'�6� �0�f�l�B���&����l��N��1��������}�D�������V�=N��U���;�9�<�
�#���������F��Y��D؊� �f�m�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h_�*���f�e�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��1��*���l�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������V��B1�L܊�d�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�����l ��h"�����3�
�`�b�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�F���
�`�e�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�����`�c�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӗ��9��h(��*���%�6�&�
�"�n�Dځ�H����g"��x)��*�����}�d�3�*����P���F��P ��U����'�:�
����������\��h��F��
�f�o����0���/����aF�N�����u�|�_�u�w�4����
����^��Q��@���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����9��h]�@���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������U��[�����u��
����2���+������Y��E��u�u�&�2�6�}��������U��N�&���������W������\F��d��Uʦ�2�4�u�0��0�F߁�����9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�(���J����CU�=��*����
����u�FϺ�����O��N�����4�u��!�%�l�>�������R��t�����
� �f�m��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��{1�� ��� �
�e�
�"�n�N߁�K����g"��x)��*�����}�d�3�*����P���F��P ��U���
�e�
� �d�d�(��Cӵ��l*��~-��0����}�e�1� �)�W���s���@��V�����!��'��8��Gہ�&����U��^�����u��
����2���+������Y��E��u�u�&�2�6�}��������l*��G1�A���0�e�3�
�a�h����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����
�:�
�:�'�o�C����֓�l ��X�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������A9��X��Eފ�
�
�
� �d�m�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����!��'��8��Gہ�&����9��h]�F���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&����\��X��G���g�0�d�a�1��A���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʲ�%�3�
�g��8�Mύ�=����z%��N�����4�u�%�&�0�>����-����l ��h_��U���
���n�w�}�����ƭ�l��h��*��d�o�����}���Y����R
��G1�����0�
��&�d�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������
F��u!��0���_�u�u�<�9�1��������V��c1��A���8�f�o����0���s���@��V�����2�7�1�g�f�}�W���5����9F������4�
�<�
�$�,�$���ƹ��^9��N��1�����_�u�w�4��������T9��S1�G���u����l�}�Wϭ�����R��^	������
�!�
�$��W���-����t/��=N��U���;�9�4�
�>�����H���$��{+��N���u�&�2�4�w�/�(���J�Г�VF��d:��9����_�u�u�>�3�Ͽ�&����A��h����������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�E��e�n�u�u�$�:����	����F��1�����u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�4��������G��h\�����o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�.����Y����V��Y1�����u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�e�w�_�w�}����Ӈ��A��E ��*���2�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�e�n�w�}�����ƭ�l��B��@���0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�e�w�]�}�W�������C9��h��U����
�����#���Q����\��XN�N���u�&�2�4�w�-��������R��N��:����_�u�u�4�0����Ӌ��v%��/��E���<�
�g�&�d�3�(���Nӯ��F�P�����}�u�u�u�w��W���7����a]ǻN��U��� �
���w�}�9���<��ƹF�N��������o��	�0���s���F�S��*����u�u����L���Y�����C1��1���o�����t�}���Y����NǻN��U���9�u�u����;���:���F�N�����o��u����>��Y���F��^ �Oʜ�u��
����2���+������Y��E��u�u�u�u�3�3�W���7ӵ��l*��~-��0����}�d�1� �)�W���s���F�T��U��������W�W���Y�ƨ�F�!��U���
���
��	�%���Hӂ��]��G��N���u�0�1�6�:�2����s���F��Z�����8�c��m���(�������]��1�<�ߊu�u�0�0�>�}�}���Y���z"�'��0���n�u�u�u�w��:���8���/��r)��N���u�u�u�1�9��>���Y�ƅ�g#��eUךU���u�u�:�!� ��?��0����v4�d��Uʥ�'�u�_�u�w�}�W���I����}F��s1��2������u�d�}�������9F�N��U���!�o�����;���:����g)��X����!�u�|�|�]�}�W���Y����\��CUװ��2�;�u�u�1�m����&�Ԣ�lU��D1�*݊�e�o�6�8�8�8�ϳ�O����'��1�����g�&�f�;��o�@���YӁ��V����U�ߊu�u�u�u��`�W��Y���F��b#��!���u�k�b�_�w�}�W����֓�z"��S�F���u�u�u�u�3�3�(���-���U��=N��U���u�:�!����J���K���F��E�����_�u�u�u�w�1�W�������XJǻN��U���0�0�u�k�6����Y���F��^ �H���'�
� �f�g�-�[���Y�����N��U���
� �f�e�'�q�W���Y����VF�	��*���f�e�6�y�w�}�W�������X��E�� ��e�%�|�_�w�}�������� T��h]����
�
�d�o�4�0����Ӌ��v%��/��E���<�
�g�&�d�3�(���N�����R��U���u�_�u�u�w�}�3��Y��ƹF�N�� �����u�k�`�W�W���Y�ƨ�]V��~*��U��f�y�u�u�w�}����&����{F�]����u�u�u�:�#�
�3���D����l�N�����4�u�_�u�w�}�W���Y����C9��\BךU���u�u�0�0�w�c����
��ƹF�N����h�u�'�
�"�n�A���U���F�
��D��u�'�
� �d�k���Y���F��RN��U���
� �f�c�4�q�W���Y����\��
P����� �f�c�%�~�W�W����֓�C��h]����
�
�g�o�4�0����Ӌ��v%��/��E���0�!�f�;��i�F���YӁ��V����U�ߊu�u�u�u��`�W��Y���F��b#��!���u�k�d�_�w�}�W����֓�z"��S�F���u�u�u�u�3�(�(���-���P��=N��U���!�8�%�}�w�}�W�������X��h�����3�
�f�
�g�W�W���Y�ƨ�F�	N�����2�
� �f�e�-�^�ԶY����lV��G��*���&�c�
�
�d�g����������r-�A���e�3�0�!�d�3�(���H�����R��U���u�_�u�u�w�}�3��Y��ƹF�N�� �����u�k�f�W�W���Y�ƨ�]V��~*��U��f�y�u�u�w�}����&����{F�X����u�:�!�8�'�u�W���Y����Z��
P��*���<�;�d�3��n�(��s���F�S��U��1�4�&�2�����L����lǑ=dךU���x�!�0�6�%�8�ϭ����R��d1�����3�!�0�&�6�8�������KǻN�����
�&�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���:����^F���&���!�
�&�
�l�}�W���Y�����Rd��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5��ԜY���F�N��U���u�4�
��1�0�K���	����U��=N��U���u�u�u�u�w�3�W���Y���F�N��U���u�3�_�u�w�}�W���Y����F�R �����0�&�_�_�w�}�ZϿ�&����A��h��ʴ�&�2�u�'�4�.�Y��s���R��R�����%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W�������]9��G��U��4�
�:�&��+�E��s���F�N�����_�u�u�u�w�}�W���Y���N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��1����|�4�1�;�#�u��������F9��W��G��4�
�:�&��+�(���P�Ƹ�V�N��U���u�u�u�u�w�}��������lV��E��I���'�
�!��%�����Iǹ��V9��1����a�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��G1�����
�
�'�2�6�.��������@H�d��Uʴ�
�0� �;�f�-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��h�� ���d�%�0�u�j�<�(���
���� T��d��U���u�u�u�0�$�W�W���Y���F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�`�3�8�f�t�������V��T��*���f�`�
�g�j�<�(���
����9��G�����u�u�u�u�w�}�W���Y�����E�����
�'�2�i�w�/�(���?����\	��^��G���d�'�2�g�b�W�W���Y���F�N��ʼ�n�_�u�u�w�}�W����ƥ�l�N��Uʰ�1�<�n�u�w�8�Ϯ�����lǑN��X���%�'�!�'����������]F��X�����x�u�u�4��8����K����T9��D��*���6�o�%�:�2�.������ƹF��R	�����u�u�u�3��-���������������h�u�d�|�#�8�}���Y���F�^�����&�u�u�d�~�)��ԜY���F�N��Uʴ�
�0� �;�e�-����DӇ��P	��C1��F؊�n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�h����H����]��X�����6�;�
� �d�h�(��DӇ��P	��C1��D��|�|�!�0�w�}�W���Y���F�N��U���'�!�'�
��/���Y����}"��v<�����g�a�0�e�%�:�E��s���F�N��U���0�1�<�n�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�u�%�%�)����&������^	�����0�&�u�x�w�}��������lU��E�����2�
�'�6�m�-����
ۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�w�l�^Ϫ����F�N��Uʼ�u�4�
�&�w�}�F�������F�N��U���u�u�4�
�2�(����	����[��G1�����9�f�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���L����lW����U���}�0�<�6�9����Lʹ��[��G1�����9�d�e�|�~�)����Y���F�N��U���u�u�%�'�#�/�(܁����F��h'��0����0�8�g�c�8�F�������l�N��U���u�u�u�0�3�4�L�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�}��������9��R	�����;�%�:�0�$�}�Z���YӇ��A��E ��*���2�4�&�2��/���	����@��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���H����[��N��U���u�u�<�u�6�����Y�����Yd��U���u�u�u�u�w�<�(�������l��PN�U���6�;�!�9�d��L���Y���F������u�u�u�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����S��D��A���;�u�:�}�2�4����&����S��G\��U���6�;�!�9�f�m�^�������9F�N��U���u�u�u�u�w�-��������C��R���������2�0�E����֓�V��\�U���u�u�u�u�w�}�������F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W��Y����V��Y1�����u�&�<�;�'�2����Y��ƹF��G1�����
�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W�������G��h[�����i�u�%�6�9�)���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�a�u�;�w�2�_ǻ�����W9��h]�L���u�u�%�6�9�)����I�����YNךU���u�u�u�u�w�}�W���	����F��1�����h�6�
����%�������l��h��*��n�u�u�u�w�}�W���YӃ����d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԶY���F��h��3����:�
�
�2��G���
������T��[���_�u�u��;���������l��h]�*���<�;�%�:�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y�ƥ�N��h��*���
�b�`�u�?�3�}���Y���F�N��U���<�
�<��%�����&���� V��S��9���
�:�
�:�'�l�A���&����l��=N��U���u�u�u�u�w�1����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y���F�^"�����'��:�
��8�(��Y����C9��Y�����e�_�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�0�3�4�L�ԜY���F��SN��N���u�0�1�%�8�8��ԶY���F��D��U���6�&�{�x�]�}�W���������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�P���Y����9F�N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�o�;���P�Ƹ�VǻN��U���u�u�u�u�e�/���A��� ��Q��Mފ�g�_�u�u�w�}�W���Y�Ɲ�r(��y-�����b�g�i�u���>�������9��d��U���u�u�u�u�w�����&����\��h\��D���2�f�m�u�j�����&����\��h\��D���
�m�
�f�]�}�W���Y���F�e��ۊ�9�
�0�:���F������� F�<�����4�9�/�'�$�o�ށ�����9��d��U���u�u�u�u�w�����&����\��h_��D���2�f�m�u�j�����&����\��h_��D���
�e�
�f�]�}�W���Y���F�^��G���2�f�c�u�j�4��������9��d��U���u�u�u�u�w�4��������U�
N����� �a�e�%�l�}�W���Y���F������
�0�
�m�n�a�W�������l ��[�����f�1�"�!�w�n�L���Y���F�N��U���0�
�0�
�`�j�K�������l ��]�����f�1�"�!�w�n�L���Y���F�N��U���c�<�
�0��e�O��Y����l��Q��E���%�n�u�u�w�}�W���Y����Q9��E��F��u�h�$�
��(�A���	��ƹF�N��U���u�u�
�
�2��O��E�ƾ�9��hY�*��_�u�u�u�w�}�W���Y����G��1����`�u�h�&�;�)��������9��d��U���u�u�u�u�w�.����	�ד�V��[�I���0�
�8�f��(�@���	��ƹF�N��U���u�u�0�
�:�n�(���&����Z�D�����b�3�
�`��o�}���Y���F�N�����d�b�'�2�d�n�W������Q��B1�C���n�u�u�u�w�}�W���YӒ��lW��h��*��`�i�u�8��l�(���O�֓�]ǻN��U���u�u�u�u�:��D�������F���*���3�
�b�
�f�W�W���Y���F�N����
�0�
�m�`�a�W���&�ޓ�F9��1��N���u�u�u�u�w�}�WϪ�	����A��V�U��!�%�a�
�"�h�C���B���F�N��U���u�8�
�f�%�:�D��Y����^��1��*��
�f�_�u�w�}�W���Y���G��^�����m�a�i�u�:��G���&����CT��N��U���u�u�u�u�#�-�A�������F���*܊� �f�m�%�l�}�W���Y����������u�u�u�;�w�;�}���Y����C��R�����u�x�u�&�>�3�������KǻN�����&�u�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��R���=�;�u�u�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��Q��M���u�=�;�u�w�}�W���Y���4��P�����:�0�
�
��i����J����[��V ��D���9�:�0�
���C���&����l��=N��U���u�u�u�u�w�/����H����lU�� N�U���0�2�d�3��e�D���B���F�N��U���u�0�0�0��3��������
F�
�����
�;�&�3��k�B���B���F�N��U���u�0�0�0��8��������R�
N�����1�/�'�&�1��B���	��ƹF�N��U���u�u�0�&�0�?��������F������a�3�
�f�b�-�_������\F��UךU���u�u�u�u�w�}��������l��h]�C��u�#�'�9� �l����A�ѓ�]ǻN��U���u�u�u�u��<�E��&���� _��R�����9�
�l�3��j�D���B���F�N��U���u�
�4�g�c�/���I�����V��A���
�f�`�%�l�}�W���Y���F���*���'�2�f�d�w�`����K����lW�� 1��N���u�u�u�u�w�}�Wϫ�����\��h��*��d�i�u�;�2�;����&����Q��G\�U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K��D��ʥ�:�0�&�u�z�}�WϮ�����N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W��PӒ��]l�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�h����H����]�R�����
� �f�`��o�JϿ�&����G9��1�\���=�;�u�u�w�}�W���Y����A��C1�����:�
�e�
���(ف�����F���*����'��:��m�(݁�&ù��U��Z����u�u�u�u�w�}�W�������G9��E1�����e�
�
�
��8�(��Y����A��C1�����:�
�e�
���(ށ�����9��d��U���u�u�u�u�w�>�(���<����G��h\�*���
�0�
�`�w�`��������A9��X��Eފ�
�
�
�
�"�n�Dց�J���F�N��U���u�6�
����%�������l��h��*��u�h�4�'�;���������R��h��*ي� �f�b�
�d�W�W���Y���F�N��*������0�:�o�A���I����lT��R�����9�
�:�
�8�-�E���K����lW��B1�Gي�f�_�u�u�w�}�W���Y�Ư�l/��r6��'���8�g�c�0�f�/���N���R��[�����:�%�g�a�e�8�F�������Q��UךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��ԶY���F��D��U���6�&�{�x�]�}�W���������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�P���Y����9F�N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�f�����P����[��N��U���u�u�u�u�4�/��������F������ �g�f�
�e�W�W���Y���F�N�����1�/�'�&�e�/���I�����R��*���:�
�
� �e�h�(��s���F�N��U���;�"�<�;�>��(���&����Z�G1��؊�e�3�
�g�d�-�_������\F��UךU���u�u�u�u�w�}�(���K����A��W�U��%��9�
�a�;�(��O����9F�N��U���u�u�u�
�6�o�D߁�����R�
N��#���
�e�3�
�e�n���Y���F�N��U���<�;�<�
�2��N��E�Ƽ�e��h\�����d�l�%�}�c�9� ���Y���9F�N��U���u�u�u�8��n�(���&����Z�G1��؊�c�3�
�e�a�-�_������\F��UךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��ԶY���F��D��U���6�&�{�x�]�}�W���������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�P���Y����9F�N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�`�;���P�Ƹ�VǻN��U���u�u�u�u��%�>�������9��P1�@���h�2�%�3��o�(��s���F�N��U���3�
����)�F�������R��S����� �f�e�%�l�}�W���Y����������u�u�u�;�w�;�}���Y����C��R�����u�x�u�&�>�3�������KǻN�����&�u�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��R���=�;�u�u�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��|�u�=�;�w�}�W���Y���F��{1��*���0��'�6�"�8�F���H¹��T9��]��Hʼ�
�!��&��)��������9��h��F��
�f�_�u�w�}�W���Y���Z*��C1�����!� �!�'��j�(ց�����^�
N��*����&�
�!�"�)����N˹��U��_����u�u�u�u�w�}�W�������l%��R1����� �0�d�`�n�/���@�����T������'�6� �2�l�B�������P��UךU���u�u�u�u�w�}��������_��S�����3�
�a�a�'�f�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠu�u�x�u�$�4�Ϯ�����F�=N��U���6�&�u�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��R��u�=�;�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��_�����e�|�u�=�9�}�W���Y���F���ي�0�
�e�f�k�}����&����T��G\�U���u�u�u�u�w�}��������l��hZ�B��u�
�4�g�c����Lù��l�N��U���u�u�u�&�;�)��������U��S�����8�`�
� �e�h�(��s���F�N��U���&�9�!�%�e�/���J�����h��@؊� �g�m�
�e�W�W���Y���F�N�����%�f�'�2�c�i�W��
����^��h��G��
�g�_�u�w�}�W���Y���G��^�����e�m�i�u�:��G���&����l��=N��U���u�u�u�u�w�0�(�������T��S�����g�3�
�a�a�-�L���Y���F���U���_�u�u�u�w�3�W���s���V��G�����_�u�u�x�w�.����	����@�CךU���'�6�&�u�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H��r�u�=�;�w�}�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�d�|�u�?�3�W���Y���F�N��*��� �!�d�'�0�i�F���DӀ��l��{:�� ��� �!�%�,�f�i�!���&����l��X�����:�`�|�_�w�}�W���Y���F��e�����
�0�
�d�c�a�W���&����g��C1�����9�
�g�
��(�E��&���F��@ ��U���n�u�u�u�w�}�W���YӖ��V��C1�����a�`�u�h�1�-����-����l+��C����b��3�
�`�k����Oӂ��]��Z����u�u�u�u�w�}�W�������l�� 1����e�u�h�3�'�%�"���6����F
��G��D����3�
�b�a�-�_������\F��UךU���u�u�u�u�w�}�(���K����A��^�U��3�%�-� ����������J9��1�����b�c�%�}�d�9� ���Y���9F�N��U���u�u�u�
�6�o�B݁�����R�
N����� ���!��1����&����e9��h\�C���}�f�1�"�#�}�E��Y���F�N��U���7�!�d�'�0�i�O���DӀ��l��{:�� ��� �!�%�,�f�i�!���&����l��_�����:�g�|�_�w�}�W���Y���F��^��*���
�d�l�i�w�%�(���5����G9��[�����g�
�
� �e�l�(��K�ƨ�D��\�N���u�u�u�u�w�}�Wϭ�����R��R	��E��i�u�0�
�:�h�(���K����CT��N��U���u�u�u�u�$�:����H����lR��N�U���
���,�"�����	����R��h��G��
�g�`�u�8�3���P���F�N��U���u�&�2�7�#�o����M����[��O��8���,� �
� �#�-���N����F9��X��G���u�:�;�:�b�t�}���Y���F�N�����d�b�'�2�c�e�W������Q��B1�AҊ�d�_�u�u�w�}�W���Y�Ƹ�C9��1����l�u�h�3�'�%�"���6����F
��G��D����3�
�b�a�-�_������\F��UךU���u�u�u�u�w�}����Mʹ��T9��Y��Hʳ�%�-� ���)�:�������T��a1��*��c�%�}�g�3�*����K��ƹF�N��U���u�u�8�
�b�����H���F��G1�� ����!��9�>�1�(��&����lT��1��]��1�"�!�u�c�f�W���Y���F�N�����`�
�0�
�f�i�K�������9��h\�G���n�u�u�u�w�}�W���YӒ��lW��h��*��l�i�u�-���;�������_��[��G݊�
� �g�d��o�B�������S��d��U���u�u�u�u�w�)���O����lR��N�U���
���,�"�����	����Q��h��G��
�g�g�u�8�3���P���F�N��U���u�!�%�d�o�/���M��� ��h��9��� �
� �!�'�$�F���/����Q��h�@���:�;�:�`�~�W�W���Y���F�N����l�'�2�a�a�}�JϷ�&����\��]����!�u�d�n�w�}�W���Y���F��u1��*���0��'�6�"�8�F�������P��S��7���
�4�0��%�>����H�ޓ�F9��\��F�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�F܁�
����O�C�����u�u�u�u�w�}�W����ԓ�9��P1�B���h�%��9��k����K�ޓ� ]ǻN��U���u�u�u�u��<�E���Hʹ��T9�� _��Hʥ��9�
�
�n�;�(��@����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�}�W��Y����]�������4�
��3�:�}�Ϫ�ӕ��G��V�����x�_�u�u�'��(���&����T��E��Oʥ�:�0�&�}�'�.����Y����`9��ZB�����y�0�<�6�9����Lʹ��l�N�����u�u�u�u�4�.�W���:����^F��=N��U���u�u�u�=�9�<�(���
�ד�@��S����u�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t�������R��C��U���%�6�;�!�;�:���P����[��N��U���u�u�u�u�w�}����*����Z�V��!���g�3�8�d�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:��؊�&�
�u�k�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W�������l ��R������&�f�3�:�o�}���Y���F�N�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�����B���F�N��U���u�;�u�3�]�}�W���Y���D����&���!�
�&�
�w�c�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�c�;���s���F�N��U���0�&�_�u�w�}�W���Y���F�V��&���8�i�u�%���܁�
����9F�N��U���u�u�u�;�w�;�}���Y���F�@��U����
�!�
�$��W���s���F�N��U���<�u�}�%�4�3��������[��G1��\���=�;�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�B�������F�N��U���u�u�0�&�]�}�W���Y���F�N������3�8�i�w�-�$���ǹ��^9��=N��U���u�u�u�u�w�3�W���s���F�N�����u�%��
�#�����Y���F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����
�&�u�h�6��#���O����lS��N��U���u�u�u�u�2�.�}���Y���F�N��U���4�
��3�:�a�W���*����9��Z1����u�u�u�u�w�}�W���Y����F�N��U���"�0�u�%���ف�
����X�N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�W���Y���F�N��U���%��
�&�w�`����-����l ��hX�U���u�u�u�u�w�}����s���F�N��U���u�u�4�
��;���Y����g9��1�����_�u�u�u�w�}�W���Y����Z ��N��U���u�u�"�0�w�-�$���Ĺ��^9��
P��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�%���.�W������l��h��*��u�u�u�u�w�}�W�������F�N��U���u�u�u�u�6��$������R��c1��B���8�c�_�u�w�}�W���Y���V��^�U���u�u�u�u� �8�W���*����9��Z1�H���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W���Y����_��N��U���u�u�u�u�w�}����*����Z�V��!���m�3�8�b�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����g9��1����h�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�VǻN��U���u�u�u�u�w�}����&����[��G1��*���e�3�8�l�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:�����3�8�l�h�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�d�1�0�F��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�F߁�
����9F�N��U���u�u�u�;�w�;�}���Y���F�@��U����
�!�d�1�0�F���G���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���;���&�u�h�4��	���&����W��N��U���u�u�u�u�2�.�}���Y���F�N��U���4�
��3�:�a�W���*����W��D��E�ߊu�u�u�u�w�}�W����ƥ�l�N��U���u�"�0�u�'��(���K����lW��
P��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�%���.�W������l��1����n�u�u�u�w�}�W���YӃ��Vl�N��U���u�u�u�u�w�<�(������F��h=����
�&�
�d�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����g9��]�����g�h�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���7����^F���&���!�a�3�8�f�f�W���Y���F�N�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�f�����K���F�N��U���u�0�1�<�l�}�W���Y�����YN��*���&�d�
�&��n�J���Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��h �����i�u�%���)�B�������9F�N��U���u�u�u�9�2�}�W���Y���F�N��U����
�&�u�j�<�(���
����U��]�U���u�u�u�u�w�}������ƹF�N��U���=�;�4�
��.�Fځ�
����[�=N��U���u�u�u�u�w�;�_���	����@��X	��*���u�%�6�|�6�9����Q����P	��h��F���
�g�h�4��2����¹��O�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���<�u�}�4��2��������F�V�����;�u�0�<�4�3�(���J����CT������!�9�d�e�~�}����Y���F�N��U���u�u�%���.�W������l��1����n�u�u�u�w�}�W���YӃ��Vl�N��U���u�u�u�u�w�<�(������F��h=����
�&�
�a�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����A�	N��U���u�u�u�u�w�}����*����Z�6��-�������u�W�W���Y�Ʃ�WF��D�U���0�1�%�:�2�.�}���Y�ԓ�l ��\�����h�&�1�9�0�>�����ι�@��R
�����;�!�9�d��n�^������]��C��F܊� �a�g�%�~�f�W���?����lU��h�I���!�
�:�<��8��������]��V�����
�#�g�a�d�}�W���������h\�� ��a�%�|�n�w�}�&���&����9��h[�*��i�u�d�u�?�3�_�������9��Q��GҊ�g�u�u�<�9�9��������_��h_�\ʰ�&�u�e�n�w�}�&���&����U��^��G��u�d�u�=�9�u����۠��U��Z��G���u�<�;�1�6�����&����lW��N�����e�n�u�u��3�ށ�����V��h��D��
�g�i�u�#�-�(���H����CT��Y
�����g�3�
�f�`�-�^�ԜY�ƞ�]��h��*���&�g�3�
�f��E��Y۴��T��V�����
�
�d�3��m�(������R��1�����0�
�
� �o�e����s���a��R_�����;�&�g�<��h����N�֓�F�F�����d�<�
� �f�n�(������R��1�����0�
�
�d�%�:�D��P���F��Y	��*���
�;�&�g�>����M����[�N��U����;�0�
�;�����K����
W��G\�����}�'�6�;�n��F���&����CT�N��R��u�9�0�_�w�}�W�������CR��Q��B܊�f�_�u�u�6�:�F�������@9��^1�*���d�g�
�g�k�}���� �ד�l ��]�*��4�1��;�2���������l��B1�Fي�f�n�u�u��3�ށ�����V��h�� ��f�
�f�i�w�}�W���YӴ��T��V�����
� �d�c��o� ���Yۉ��P	��]��*���d�`�
�g�g�}�W��PӃ��VFǻN��U���0�
�8�g��(�F��&����F�e��ۊ�9�
�;�&�e�0����&����Q��G\��H���4�2�d�4�;�2����&�ד�V��V����6�'�,�d�9�)�ށ�����9��UךU���4�2�d�4�;�2����&����Z9��h_�@���u�h�}�4�0�l��������9��Q��@���%�u�;�u�6�/�(ށ�����U��Y�����_�u�u�4�0�l�������� 9��hV�*��i�u�!�%��(�O���	�ƭ�WF��G1�*���m�m�%�|�]�}�W����ד�_
��Y��@���
�l�c�%�w�`�U���������R�����'�2�a�d�w�}��������EU��N�����e�n�u�u��3�ށ�����V��h��F��
�g�i�u�f�}����Q����@��hZ�����d�l�h�4��2����������RN��W�ߊu�u�4�2�f�<��������lW��1��U��}�4�2�g�6�1����&¹��U��[�����;�u�4�2�f�<��������U��W�����_�u�u�4�0�l��������lW��B1�Lߊ�g�i�u�d�w�5��������U��]�����u�%�6�;�#�1�Bہ�PӃ��VF�UךU���4�2�d�4�;�'����K����
T��G\��H���4�2�d�4�;�2����&����^��N��ʴ�
�:�&�
�!��^�ԜY�ƞ�]��h��*���:�
�
�d�1��G���	���l�N��Uʥ�l�
�d�3��n�(������	��T��Lي�d�3�
�d��o�G���Y�����RNךU���u�u�0�
�:�i�(���@�ԓ� ]ǻN�����d�4�9�/�%�.�E�������_��N�U���u�u�u�%�n��(���H����CT��_��]���6�;�l�
��(�F��&���F�_��U���0�_�u�u�w�}��������U��Z����u�u��;�2��������� 9��hW�*��i�u�d�u�?�3�_���&����U��Z��F��4�
�:�&��+�C��Y����D��d��Uʇ�;�0�
�9��8����&����
U��G\��H���w�"�0�u�'�����&¹��T9��\��U���6�;�!�9�d�m�W�������l�N�����
�9�
�0�8��(���J����CT�
N��Wʢ�0�u�%��$�1�(ہ�����_������!�9�f�e�w�1����[���F��Y	��*���
�0�:�
�"�l�@؁�K���4��P�����:�0�
�
�"�l�N؁�KӞ����T�����d�d�n�u�w�����&����U��]�����h�&�1�9�0�>�����ο�Z ��E�� �&�2�0�}�6��(���H����CU�C�����0�}�;�<�9�9�P���_Ӓ��lT��Q��A���%�}�d�d�3�*����P���l�N�����
�
�
� �o�i����Dӕ��l
��^�����'�&�<�!�%�:�ǫ�
����WN��Y1��C���
�d�
�f�{�2��������]��Y��R��s�!�%�c��(�O���	����W��X����|�|�n�u�w�����&����\��h_�� ��c�%�u�h�u�� ���Y۴��T��a1�����m�
�g�h�%��F���&����CT�R��U��n�u�u��9�8�(���&����lW��1��*��
�f�i�u�w�}�W���+����9��[1�����
� �m�c�'�}����Q����\��1��*���m�a�%�}�~�`�P���Y����l�N��Uʧ�#�
� �m�e�-�L���YӴ��T��V�����
�
�
� �f�h�(��E��ƹF�N�����g�4�9�:�2����Mƹ����YN�����;�l�
�
�"�l�E܁�K���F�G�����_�u�u�u�w�8�F���&����l��=N��U���2�g�4�9�8�8�(ށ�����l ��Y�*��i�u��;�2���������l��E��F��u�:�u�%�4�3����H���9F�<�����4�9�:�0������&����^��G\��H���4�2�g�4�;�2����&����lW��1��U���u�%�6�;�#�1�F��B���4��P�����:�0�
�
�"�o�Eށ�K���W�@��U¥��&�9�
��j����M����F��h�����#�
�|�0�$�}�G��Y����R��1�����0�
�
� �d�m�(��E���F��R �����&�9�
�
�2��F��DӇ��P	��C1��G��u�9�0�w�u�W�W�������l��h�����
�a�`�%�w�`�U�������4��P��#���3�
�a�f�'�}�W���&����U��G\�����u�e�n�_�w�}�ZϿ�&������^	�����0�&�u�x�w�}��������@��Y1�����u�'�6�&��-�����ƭ�l��h�����
�!�
�&��q�����ƭ�l��h�����
�!�`�3�:�l�[ϻ�����W9��h]�L���|�u�u�7�0�3�W���Y����UF� ��]´�
�:�&�
�8�4�(���Y����G��G�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�W���Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�4�
�<��.����&����l ��h_�U���u�:�}�0�>�>��������
9��S�����;�!�9�d�g�t�^������F�N��U���4�
�:�0�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����S��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C�����9�u�&�<�9�-����
���9F������
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9��=N��U���<�_�u�u�w�}�������R��X ��*���<�
�u�u�'�.����PӇ��N��h�����:�<�
�u�w�-��������`2��C_�����|�|�!�0�w�}�W���Y�����^
��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}���������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����V�������%�:�0�&�w�p�W�������R��V�����'�6�o�%�8�8�ǿ�&���R��^	������
�!�`�1�0�F������\��Q��A���%�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��Dߊ�&�
�a�u�9�}��������\��Q��A���%�u�u�%�4�3����H���O��_�����u�u�u�u�w�-���� ���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�'�4�,�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��8����IӇ��Z��G�����u�x�u�u�6������֓�@��Y1�����u�'�6�&��-�������T9��R��!���d�
�&�
�c�}��������F9��W��G���'�
�!��%�����Iǹ��V9��1����a�u�%�'�#�/�(߁����F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O��Y
�����0�<�6�;��(�D��&�����T�����d�e�|�|�#�8�W���Y���F������'�
�u�h�6�/��������\��Z��*���
�
�0�
�a�f�W���Y����_��=N��U���u�u�u�%�%�)����Y����C9��C��*ڊ�'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����F��N�����u�'�6�&�y�p�}���Y����V��Y1�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�h����H����K��X �����a�l�%�y�6�/��������\��Z��*���
�0�
�b�{�<�(�������l��PGךU���0�<�_�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\ʴ�1�;�!�}�/�)��������_��N�����:�&�
�#��t�^������F�N��U���4�
�0� �9�l�K�������l ��h"����a�g�0�d�%�:�E��s���F�R��U���u�u�u�u�w�<�(�������Z�V�����;�d�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��C��*���&�<�;�%�8�8����T�����E�����
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	���&����R�R�����
� �f�`��o�W���0����r4��R��G���0�e�'�2�e�n�W�������]9��G��\���u�7�2�;�w�}�W��������T�����2�6�d�h�6���������C9��Y�����6�d�h�4��4�(�������@��h��*��u�;�u�:��8��������lU��1��U���%�6�;�!�;�l�G���PӒ��]FǻN��U���u�u�%�'�#�/�(���DӅ��z(��o/�����
�f�
�
��8�(��B���F����ߊu�u�u�u�w�}��������F������'�
�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��R����4�&�2�u�%�>���T���F��h�� ���f�4�&�2��/���	����@��G1��Yʴ�
�<�
�&�&��(���L����lW�������1�3�
�a�n�-�[Ͻ�&����k'��C��*��
�
�
�0��e�[Ͽ�&����A��h���ߊu�u�0�<�]�}�W���Y���N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��1����|�4�1�;�#�u��������F9��W��G��4�
�:�&��+�(���P�Ƹ�V�N��U���u�u�4�
�2�(���E�Ư�l/��r6��'���8�g�a�0�f�/���O���F�N�����u�u�u�u�w�}��������lU�
N��*��� �;�f�%�2�f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����E�����u�&�<�;�'�2����Y��ƹF��G1�����
�
�&�<�9�-����Y����V��V�����%�&�2�6�2��#���Hƹ��^9��N�����;�
� �f�b��E�������v>��e����c�0�e�'�0�o�E���	����F��1�����u�u�7�2�9�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��[�����a�u�;�u�8�u��������U��[�����u�%�6�;�#�1�F��P����[��=N��U���u�u�u�%�%�)����Y����_9��s+��'���'�
�f�
������M��ƹF�N�����_�u�u�u�w�}�W�������]9��S�����!�'�
�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h�� ���`�4�&�2�w�/����W���F�V�����;�`�4�&�0�����CӖ��P�������4�
�<�
�$�,�$����ӓ�@��B�����:�1�3�
�c�d�������w#��e<�����f�
�
�
�2��N������G��h[�����_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C_�����d�|�4�1�9�)�_�������l ��Z�*��h�4�
�:�$��ށ�P���G��d��U���u�u�u�4��8����L���P
��y*��4���0�8�g�c�2�l����K����F�N�����u�u�u�u�w�}�WϿ�&����A��R�����0� �;�`�'�8�L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����1�d�`�4�$�:�W�������K��N�����<�
�1�
�d���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����J���N��h�����#�
�u�u�'��(���Q�ƨ�D��V��N���u�0�1�%�8�8��Զs���K��G1�����1�d�f�4�$�:�W�������K��N�����<�
�1�
�a���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����O���N��h�����#�
�u�u�'��(���Q�ƨ�D��W��N���u�0�1�%�8�8��Զs���K��G1�����1�d�`�4�$�:�W�������K��N�����<�
�1�
�o���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����A���N��h�����#�
�u�u�'��(���Q����\��XN�\��u�u�0�1�'�2����s���F������7�1�g�b�6�.��������@H�d��Uʴ�
�<�
�1��m�(�������A	��N�����&�4�
��1�0�}���Y����]l�N��U���u�u�u�4��4�(���&����[�V�����
�#�
�u�w�-�4���
������Y��D���n�u�u�0�3�-����
��ƓF�C�����2�7�1�g�g�}����Ӗ��P��N����u�%�&�2�5�9�E��&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����W��R��]���6�;�!�9�f�l�JϿ�&����@�
�����d�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��l�NϿ�
����C��R��U���u�u�4�
�>�����H�ߓ�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��^�I���4�
�:�&��+�(���Y����`9��ZF����!�u�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�E��Y����T��E�����x�_�u�u�'�.��������9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�D���h�}�%�6�9�)����H����C9��h��]���:�;�:�f�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����H����@��YN�����&�u�x�u�w�<�(���&����W��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��a�i�u�4��2����¹��F��h-�����a�1�"�!�w�t�L���YӃ����T��N�ߠu�u�x�u�'�.��������F��D��U���6�&�{�x�]�}�W���
����W��]�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����g�f�u�h��-��������lW���6���&�}�u�:�9�2�B���s���V��G�����_�_�u�u�z�<�(���&����S��V�����'�6�&�{�z�W�W���	����l��h\�*���<�;�%�:�w�}����
�έ�l%��Q�����u�0�<�_�w�}�W���Y���F��h��*���
�`�u�h��-��������lW���6���&�}�g�1� �)�W��P���F��SN�����&�_�_�u�w�p��������W9��N�����u�'�6�&�y�p�}���Y����Z��S
��Bۊ�&�<�;�%�8�}�W�������R��d1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�b�u�j�u��������EW��S�����
�&�}�f�3�*����J����F�R �����0�&�_�_�w�}�ZϿ�&����Q��Y�U���<�;�%�:�2�.�W��Y����C9��P1����a�
�&�<�9�-����Y����V��V�����&�$��
�#�h����H����K��X �����a�l�%�|�w�}�������F�N��U���u�%�&�2�5�9�E��Y�����T�����2�6�d�h�6�����
����g9��[�����a�u�;�u�2�4����&����S��G\��U���6�;�!�9�f�m�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��Y�����;�%�:�u�w�/����Q����`9��ZGךU���0�<�_�u�w�}�W���Y���R��^	�����m�u�h�}�'�>�����ד�[��G1��*���}�a�1�"�#�}�C���s���V��G�����_�_�u�u�z�<�(���&���� U��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��]�����;�%�:�u�w�/����Q����`9��ZGךU���0�<�_�u�w�}�W���Y���R��^	�����f�i�u�4������Iӂ��]��G��U���6�;�!�9�f�l�L���YӃ����T��N�ߠu�u�x�u�'�.��������R��P �����&�{�x�_�w�}��������lP��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��C���h�}�%�6�9�)����H����C9��h��]���:�;�:�c�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����HӇ��Z��G�����u�x�u�u�6���������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��hV�I���4�
�:�&��+�(���Y����`9��ZF����!�u�|�n�w�}����	����@��=d��U���u�%�&�2�4�8�(���
����U��N�����u�'�6�&�y�p�}���Y����Z��D��&���!�e�3�8�n�<����&����\��E�����%�&�2�7�3�l�D�ԜY�Ʈ�T��N��U���<�u�4�
�>�����O����[��=N��U���u�u�u�%�$�:����&����GW��Q��L��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}��������V��c1��Dڊ�&�
�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�>����-����9��Z1�U���<�;�%�:�2�.�W��Y����C9��P1������&�d�
�$��G���
����C��T�����&�}�%�&�0�?���L���F��P��U���u�u�<�u�6���������O��_�����u�u�u�u�w�-��������`2��C_�����d�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����Z��D��&���!�d�3�8�f�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��C_�����d�u�&�<�9�-����
���9F������6�0�
��$�l�(���&�ד�@��Y1�����u�'�6�&��-��������Q�N�����;�u�u�u�w�4�Wǿ�&����Q��^�U���;�_�u�u�w�}�W���	����l��F1��*���g�3�8�d�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h��*���$��
�!�e�;���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��F1��*���f�3�8�d�w�.����	����@�CךU���%�&�2�6�2��#���H����^9��h�����%�:�u�u�%�>����	����l��h\�\���u�7�2�;�w�}�W�������C9��P1����l�u�=�;�]�}�W���Y���R��^	������
�!�f�1�0�F���DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����<�
�&�$����������F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��^	������
�!�a�1�0�F���
������T��[���_�u�u�%�$�:����&����GW��Q��Dي�&�<�;�%�8�}�W�������R��^	�����b�|�u�u�5�:����Y����������7�1�g�d�w�5��ԜY���F�N��*���
�&�$���)�C�������[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����l ��h_�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���
�&�$���)�B�������R��P �����&�{�x�_�w�}��������B9��h��@���8�d�
�&�>�3����Y�Ƽ�\��DF��*���
�1�
�m�~�}�Wϼ���ƹF�N�����%�&�2�7�3�o�@������F�N��U���4�
�<�
�$�,�$����ӓ�@��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����
����g9��[�����a�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�<�
�$�,�$���¹��^9��V�����'�6�&�{�z�W�W���	����l��F1��*���
�&�
�
�$�4��������C��R�����<�
�1�
�d�W�W�������F�N�����4�
�<�
�3��D������F�N��U���4�
�<�
�$�,�$���¹��^9��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��Q��E��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���݁�
����R��P �����&�{�x�_�w�}��������B9��h��*���
�
�&�<�9�-����Y����V��V�����1�
�d�d�]�}�W������F�N��U´�
�<�
�1��l�F������F�N��U���4�
�<�
�$�,�$�������^9��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��Q��D��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���܁�
����R��P �����&�{�x�_�w�}��������B9��h��*���
�
�&�<�9�-����Y����V��V�����1�
�d�l�]�}�W������F�N��U´�
�<�
�1��l�N������F�N��U���4�
�<�
�$�,�$�������^9��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��Q��G��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���ہ�
����R��P �����&�{�x�_�w�}��������B9��h��*���
�
�&�<�9�-����Y����V��V�����1�
�d�b�]�}�W������F�N��U´�
�<�
�1��l�@������F�N��U���4�
�<�
�$�,�$���ǹ��^9��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��Q��F��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���ځ�
����R��P �����&�{�x�_�w�}��������B9��h��*���
�
�&�<�9�-����Y����V��V�����1�
�d�a�]�}�W������F�N��U´�
�<�
�1��l�C������F�N��U���4�
�<�
�$�,�$���ƹ��^9��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��Q��A��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���ف�
����R��P �����&�{�x�_�w�}��������B9��h��*���
�
�&�<�9�-����Y����V��V�����1�
�d�g�]�}�W������F�N��U´�
�<�
�1��l�E������F�N��U���4�
�<�
�$�,�$���Ź��^9��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��Q��@��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���؁�
����R��P �����&�{�x�_�w�}��������B9��h��*���
�
�&�<�9�-����Y����V��V�����1�
�l�_�w�}����s���F�^�����<�
�1�
�n�}����s���F�N�����<�
�&�$���؁�
����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����U��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�V�����&�$��
�#�����Y����T��E�����x�_�u�u�'�.��������l��h��*݊�&�<�;�%�8�}�W�������R��^	�����d�_�u�u�2�4�}���Y���Z �V�����1�
�d�u�?�3�}���Y���F�V�����&�$��
�#�����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�<�
�&�&��(���&����F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��^	������
�!�
�$��W�������A	��D�X�ߊu�u�%�&�0�>����-����l ��hV�����;�%�:�u�w�/����Q����Z��S
��F���u�u�7�2�9�}�W���Yӏ����D�����d�`�u�=�9�W�W���Y���F��h��*���$��
�!��.�(���DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����<�
�&�$���ց�
����[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���Y�ƭ�A9��h(��*���%�g�a�e�2�m����O�ӓ�F���*���<�
�0�!�%�/����Q����V��Z��Eފ� �f�l�
�c�q�E���s�����h��3����:�
�e���(ށ�����
9��R�����9�2�6�#�4�2�_���������C��D���
�4�2�
�9������ԓ�F9��\��F���u�;�<�;�3�<����&����	��h\�*ڊ�
�
� �f�g��F���s���R��[�����:�%�g�a�e�8�G�������U��N�U���u�u�u�6���2���+����lT��h��*���
�a�u�=�9�u�����ԓ�F9��]��G��u�u�d�|�2�.�W���Y�����h��3����:�
�e���(߁�����9��d��Uʴ�'�9�
�:��2���M�ԓ�lV��h��F��
�f�i�u�w�}�W�������G9��E1�����e�
�
�
��(�D��&����[����*���
� �f�b��o�G���Y�����RNךU���u�u�9����%�������9��1����f�_�u�u�%���������C9��1�����f�3�
�c�n�-�W��s���F�T��;�����0�8�e�i��������U��_��]���
�8�g�3��i�D���Q���A��N�����u�u�u�u�6�/��������\��Z��*���
�
� �f�d��D�ԜY�ƭ�A9��h(��*���%�g�a�g�2�m�B���&����l��S��U���u�u�4�'�;���������R��h��*���f�e�
�d� �8�Wǭ�����9��h]�F���}�|�h�r�p�}����s���F�V�����:�
�:�%�e�i�E���I�Г�V��Z�U���4�'�9�
�8�����K�ғ�l��h��F��
�f�i�u�w�}�W�������w#��e<�����f�
�
�
�2��C������@��C�����a�d�%�}�~�`�P���Y����l�N��Uʴ�'�9�
�:��2���M�֓�lV��B1�Eߊ�d�_�u�u�%���������C9��1�����d�3�
�c�b�-�W��s���F�V�����:�
�:�%�e�i�G���H���� P��h����u�&�9�!�'����A����V�
N��R���9�0�_�u�w�}�W���&����\��X��G���g�0�d�'�0�o�B�ԜY�ƭ�A9��h(��*���%�g�a�g�2�l�E���&����l��S��U���u�u�4�'�;���������R��h��*���f�e�
�g� �8�Wǭ�����l ��Z�*��e�u�u�d�~�8����Y���F��[1��1����!�'�
�d��(ށ�����]ǻN�����!��'��8��Gہ�&���� 9��h]�D���u�h�_�u�w�}�W���0����r4��R��G���0�d�'�2�e�k� ���Yە��l��1��*��f�%�}�|�j�z�P������F�N�����9�
�:�
�8�-�E���K����lT��B1�Cي�f�_�u�u�%���������C9��1�����a�3�
�c�n�-�W��s���F�T��;�����0�8�e�k��������
Q��_��]���
�8�
� �d�j�(��I���W����ߊu�u�u�u�%���������C9��1�����3�
�c�l�'�f�W�������G9��E1�����e�
�
�
�����AĹ��Z�=N��U���u�9��������&����V9��E��G��"�0�u�&�;�)�݁����� 9��^��H��r�u�9�0�]�}�W���Y����_��X�����g�a�g�0�f�i����O�ߓ� ]ǻN�����-���!��8����6����F��1��*��c�%�u�h��0�(��&���� S��G]�����%�6�;�!�;�l�F��Y����\	��O)��:����0�!�'������&����lT�� 1��U��}�8�
�f��8�(��HӞ����T�����d�d�n�u�w�?����>����G9��R�����
�$�4�
��(�E��&���F��[�� ��l�
�g�-�%�<�(���
����9��d��Uʷ�8�'�0�
�"�l�N܁�K�����_�� ��m�
�g�:�w�/����@Ĺ��^	��V ��D���
�m�f�%�~�W�W�������VR��S�����
�d�3�
�n�o����D�΢�D��Y��*ي� �g�e�
�d�<�Ϻ�����l	��D1�����l�`�%�|�]�}�W�������9��Z�����g�3�
�d�f�-�W��Q����Z��^��*���f�m�
�f�6�9��������]��1��*��a�%�|�_�w�}��������W��E	��*��� �g�e�
�e�a�Wǭ�����l��h]�Cʴ�1�;�"�<�9�4�(݁�����
V�=N��U���0�2�l�
�2�2����¹��lW��1��U��}�0�&�2�5�)�F���&����l��V �����!�1�:�0���F���&����l��d��Uʷ�8�'�0�b�3�0����&����lW��1��U��}�0�&�2�5�)����J����R��S�����:�0�
�
��(�F��&���9F������l�
�d�3��e�N���Y���Q��E	��B���8�'�4�
�f�;�(��J����K	��V�����
�#�
�|�]�}�W�������9��Q��L���%�u�h�}�%�8���&����A��h�� ��c�
�g�-�%�<�(���
����9��d��Uʷ�8�'�0�l�>����N����Z������
�:�
�d�1��@���	�ƣ�4��P�����:�0�
�
�8��F���&����l��d��Uʷ�8�'�0�l�>�;�(��@����[�T�����;�!�<�3��h�@���Y����R��1�����0�
�
�:�����A����]ǻN�����2�
� �d�n��E��Yے��9��h_�D���u�'�7�8�%�8�@�������]9��Q��L���%�|�_�u�w�/����&�ד�F9��X��G��u�;�"�<�9�4�(ށ�����9�������!�1�/�'�$�m����¹��lW��1��\�ߊu�u�'�0�0��E���&����l��S�����<�;�<�
��8�(��IӉ��C9��C1�����g�m�%�|�]�}�W�������ZU��B1�Bߊ�g�i�u�;� �4����&����lT��1��U���%�;�!�<��(�E��&���9F������
�a�3�
�f�i����D�΢�D��Y��*ފ� �f�m�
�d�2�W�������l ��_�*��n�u�u�7�:�/��������P��N�U»�"�<�;�<��8�(��IӉ��W��C�����&�e�;�!�>�;�(��H����l�N�����0�<�<�
�"�o�Aہ�K�����R�����
�0�
�l�f�2�W�������lW��R	��L��n�u�u�7�:�/��������lT��1��U��}�;�0�3�8��(���K����CT��EN�����:�
�
� �e�d�(��B�����R��*���f�3�
�e�b�-�W��Q����A ��@1�����e�e�%�u�%�2��������U��V�����_�u�u�'�2�:�(���M���� W��h�I��� �1�'�9� �i����H�ߓ�F�������"�a�3�
�f�h����s���Q��E	�����3�
�l�l�'�}�J�������_	��Q��L���%�u�'�:�2�;��������9��UךU���4�'�
�
�"�o�Fف�K�����h_�*���
�e�g�4�3�)���&����
W��G\����u�4�'�
��l����N�֓�F�F�����%�g�3�
�a�o�����Ƹ�CQ��B1�Gފ�g�n�u�u�4�/��������U��h�I���&�9�!�%�f�;�(��I����R��C��*���d�d�
�g�l�}�WϽ�����l��h�����b�d�%�u�j�u��������P��N��U���
�g�
� �f�j�(��B�����E��*���
�
� �d�`��E��Yے�� 9��h_�D���u�'�!�%�`����J����]ǻN�����
�
� �f�n��E��Yے��lW��h��*��l�4�1�!�'�d�(���J����CT�=N��U���'�
� �g�d��E��Yے��lW��h��G��
�f�4�1�#�-�@ځ�����9��UךU���
�&�<�;�f�;�(��&���F��h��#���!�d�m�'�0�n�B��Y����l��^	�����f�
�e�i�w����� ����T��E��F��n�u�u�1�;�)��������ZW��B1�E܊�g�i�u�1�;�)��������U�� V�����'�&�9�!�'�o����A�ד�O��N�����!�1�:�0���(���H����CT�
N�����0�
�;�&�%�:�D��Y����V
��Z�*���d�e�
�g�l�}�WϺ�����l	��D1�����b�f�%�u�j�W�W���Y�ƞ�]��h��*���&�g�8�-�>����N˹����YN�����2�l�
�d�1��@���	����[�I�����u�u�u�u�w�-�Nف�H����lU��UךU���0�0�0�
�9�.�E���&����l��S��U���u�u�%�a��l����@�ߓ�F��R �����,�d�3�
�n�k����P���A�R��U���u�u�u��9�8�(���&����lS��B1�G܊�g�_�u�u�2�8��������l ��_�*��i�u�u�u�w�}���&�ԓ�F9��V��Gʢ�0�u�6�'�.�o����I�ӓ�N��S��D���0�&�u�u�w�}�Wό�����R
��X ��*܊� �f�e�
�e�W�W�������W9��R�� ��d�
�f�i�w�}�W���YӴ��T��V�����
�
� �
��(�F��&����[�������l�
�
� �f�e�(��I���W����ߊu�u�u�u��k����&����l��=N��U���0�0�
�0�8��(���&�ד�F9��_��G��u�!�%�c��8�(��MӇ����R��*���:�
�
�:��(�F��&���9F�
�����
�0�:�
��2�(�������9��R��]���
�g�'�2�d�l�W���Y����G��M�����!�3�
�l�a�-�^�ԜY�ƨ�_��S1�����d�3�
�b�c�-�W��s���F�e��ۊ�9�
�;�&�e�4�(���&������YN�����
�
�d�3��j�G���Q���A��N�����u�u�u�u��3�ށ�����A	��1��*���
�m�f�_�w�}��������A	��1�����
�m�`�%�w�`�_�������I��D1�����b�a�%�u�8�}��������EW��UךU���0�0�0�
�2�2�(݁�����9��R��]���;�<�
� �e�i�(������\��V��*���g�a�
�g�l�}�WϺ�����l��X��*���g�f�
�f�k�}�W���Y����R��1�����0�
�
� �e�o�(��������E��*���g�d�
�g�g�}�W��PӃ��VFǻN��U���4�2�d�4�;�'����M����_��h����u�0�0�0��8����&����W��G]��H�ߊu�u�u�u�6�:�F�������@9��Q��D���%�u�=�;��<����&����_��G\��\��r�r�u�9�2�W�W���Y�ƞ�]��h��*���:�
�
� �d�l�(��s���W��C�����&�3�
�`�`�-�W��s���F�e��ۊ�9�
�;�&�e�4����L�Փ� F��R �����,�d�<�3��n�B���Q���A��N�����u�u�u�u��3�ށ�����A	��1�����`�l�%�n�w�}��������V��h ��*���d�f�
�g�k�}��������V��h��*��a�-�'�4��2����¹��l�N�����;�
� �f�b��E��Y���D��F��*����'��:������I���R��X ��*���
�|�0�&�w�m�L���YӃ��l0��h��A���%�u�h�&�3�1��������AN��D�����8�
�c�3��e�(��Y�ƹ�@��R
�����;�!�9�d��m�^��Y����K��h��F���%�u�h�&�3�1��������AN��D�����8�
�
� �d�i����Rӓ��Z��SF��*���&�
�#�g��l�^�ԜY�Ʃ�C9��G1��D���
�b�
�a�k�}����/�ד�F9��1��]��1�"�!�u�e�f�W�������^��h��F���%�u�h�<�2��(���J�ޓ�N��
�����`�|�_�u�w�%�(�������r��[��*��� �
�b�d�1��E���	���l�N��Uʥ��9�
�c�%�:�D��Y����N��G1�*���g�c�
�g�g�}�W��PӃ��VFǻN��U���-�
��-�"���������R
��hW�����
�g�b�%�l�}�Wϸ�	����K)��h/�����0��9�0�n��(���K����CT�
N�����2�6�#�6�8�u��������C9��Y����
�|�x� �$�:����&����lW��E��F��|�n�u�u�1�-�6���6����Q��B��#���0�l�
�
�"�o�Oہ�J���9F�N��U���4�g�a�
�"�o�B߁�Jӑ��]F��Z��B���
�f�g�%��t�J���^�Ʃ�@�N��U���3�%����)�6�������e��R1�*��� �g�b�
�e�W�W�������`��C1�����!�
�4� ��d����&����l��S�����:�<�
�0�#�/��������R��X ��*���a�e�u�u�9�4����	����9��h��G���
�f�|�_�w�}��������V��W��#���
�`�f�%�w�`��������l��C�� ���2�0�}�%�4�3����Kƹ��K��Y�����3�%�;�1��8���I����F9��^��D���_�u�u�-��2��������9��Q��@���%�u�h�&�3�1��������AN��D�����%�6�;�!�;�o�(���Tӓ��Z��SF�����1�
�0�8�b�k�!���&����l��UךU���u�u�-�
�8�8����&����e9��h\�L���u�h�&�1�;�:��������A��M�����1�%��9��l����M����T��UװU���u�u�3�%�9�9�(�������l0��B1�Eڊ�d�i�u�!��2����������^�����0�}�
�4�e�l�(���&����J��G����u�-�
�0�:��Cہ�&����W��G]��H�ߊu�u�u�u��<�E��&����U��X�����=�;�}�0��0�Cׁ�����9��^��H��r�u�9�0�]�}�W���Y����G��1��*��b�%�n�u�w�;����,����F��B�����d�a��3��j�A���Y����^��1��*��g�%�}�g�z�l��������l�N����� ���!��1����&����e9��h\�C���u�h�'��c�;�(��A����9F���*����,� �
�"�)����H�ғ�l ��Y�*��i�u�!�
�8�4�(�������V��RF�����0�}�!�
�8�4�(�������Z��SF����� ���!��1����&����e9��h\�C���|��&�2�2�u����4����|��z�����
�g�
�
�"�o�Gف�H���S��UךU���-�
���.�(�(�������lW��h8�� ��d�
�e�i�w�0�(�������T��F�U���u�:�;�:�g�f�W�������~3��N!��*���!�%�,�d�`�����N�Г�F���*ߊ� �g�l�
�e�W�W�������f*��x��8���<�9�
�g�����HŹ��Z�D�����6�#�6�:��8��������]��D�����6�#�6�:��4��������~3��N!��*���!�%�,�d�`�����N�Г�O������3�%�-� ����������J9�� 1�����b�c�%�|�~�}�@���s���K�P�����g�
�0�4�$�:�W�������K��N�����3�
�g�
�2�<����&����\��E�����%�&�4�!�w�-��������`2��C_�����y�4�
�0�w�-��������`2��CY�����y�4�
�<��.����&����U��B�����2�6�0�
��.�D������R��^	������
�!�
�$��[Ͽ�&����P��h=�����3�8�a�u�'�.��������l��h��*���u�u�7�2�9�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����N��G1�����9�2�6�d�j�<�(���&����l5��D�����e�u�;�u�8�u��������F��h�����:�<�
�|�~�2�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���Ĺ��^9����]���6�;�!�9�0�>�F������T9��R��!���g�3�8�d�w�/�_�������l
��^��U���%�&�2�6�2��#���J����lT�X�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�8�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��EN�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�`�|�~�)����Y���F�N����� �f�e�6�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��G1��*��
�0�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=d��Uʲ�%�3�
�g��m�K�������l��_��N���u�2�%�3��o�(��E�ƥ�l��h��*��_�u�u�x�0�-����KŹ����^	�����0�&�u�x�w�}��������9��h�����%�:�u�u�%�>����	����A�V�����&�$��
�#�����UӇ��P�V�����&�$��
�#�����UӇ��@��T��*���&�g�3�8�f�}��������B9��h��*���
�y�4�
�>�����*����9��Z1�U���&�2�6�0��	��������F��h��*���$��
�!��.�(���Y����V��=N��U���u�3�}�}�'�>��������lW������4�1�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��CF�����4�!�h�4��2��������O���]���6�;�!�9�0�>�F������T9��R��!���b�3�8�c�w�/�_�������l
��^��U���%�&�2�6�2��#���K����lW�X�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�8�}��������_	��T1�Hʴ�
�<�
�&�&��(���&���� O��EN�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�a�u�%�u��������\��h_��U���&�2�6�0��	��������O����ߊu�u�u�u�w�}��������l��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�2�'�;�(��&���F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�}�WϹ�	���� T��G^��Hʼ�
�0�
�0�6�m�}���Y����U��X��D��u�;�'�3�:�%�D�ԜY�ƥ�l��t��*��� �!�'�
�`��G���&����l��S�����:�<�
�0�#�/�����Υ�l��t��*��� �!�'�
�`��(���J����CW�N�����}�
�4�g�$�l�(���&����O��N�����!��&�
�#�(����&����W��B1�M؊�f�i�u�u�w�}�WϷ�&����R��d�����0�d�d�d��(�D��&����[����*���c�
� �f�`��E��Y���O��[�����u�u�u��4�����*����G��h_�*ي� �f�`�
�d�W�W���5����p��h=�� ���'�
�b�
�e�;�(��@����[�N��U���<�
�!��$���������^��1����l�u�=�;��8�(���K���� R��h�E���u�d�|�0�$�}�W���Y����9��h-�����'�6� �0�f�l�B���&����l��=N��U���6�
�4�0��/��������lW��B1�Dڊ�f�i�u�u�w�}�WϷ�&����R��d�����0�d�m�m�1��E���	�ƻ�V�C��Lӊ� �f�c�
�e�m�W���H����_��=N��U���u��6�
�6�8�$�������lW��h��F��
�f�_�u�w���������G��C��*��
�
� �f�d��D��Y���F������4�0��'�4�(���L�ޓ�F9��Z��Gʢ�0�u�&�9�#�-�N���&����l��G��U��|�0�&�u�w�}�W�������l%��R1����� �0�d�d�f�;�(��I����9F������4�0��'�4�(���H�Փ�F9��X��F��u�u�u�u�w�4�(���:����`��T����m�m�3�
�e�h�������@��C��D���
�f�e�%��t�J���^�Ʃ�@�N��U���<�
�!��$���������Q��1��*��e�%�n�u�w�4�(���:����`��T����d�`�3�
�c�j����D���F�N��*����&�
�!�"�)����N˹��A��_�U���;�}�0�
�:����N¹��V�
N��R���9�0�_�u�w�}�W�������@��C�����
�b�
�d�%�:�C��B�����T������'�6� �2�l�F���&����l��S��U���u�u�<�
�#���������F��Y��Dڊ� �f�`�
�e�*����
����^��h��*��c�e�u�u�f�t����Y���F������4�0��'�4�(���L�ޓ�F9��Z��G�ߊu�u��6��<��������A�� V��*���f�l�
�f�k�}�W���Y����9��h-�����'�6� �0�f�h�O���&����l��@��U¡�%�l�
� �d�k�(��I���W����ߊu�u�u�u��>�(�������F��E��BҊ� �f�l�
�d�W�W���5����p��h=�� ���'�
�b�
��(�D��&���FǻN��U����6�
�4�2���������^��h��F���
�d�"�0�w�.����	�ߓ�F9��Z��G��u�u�d�|�2�.�W���Y�����T������'�6� �2�l�O�������
V��UךU����6�
�4�2���������^��h��F��
�f�i�u�w�}�W�������l%��R1����� �0�d�d�f����Lʹ����YN�����8�c�
� �d�h�(��I���W����ߊu�u�u�u��>�(�������F��E��BҊ�
� �f�l��n�}���Y���Z*��C1�����!� �!�'��j�(ׁ�����9��R�����9�2�6�#�4�2�_�������Z��SF����
� �f�a��i�[��P��ƹF��{1��*���0��'�6�"�8�F���@���� R��h�I���u�u�u�u�>�����
����A��B��D���m�3�
�g�c�-�W����ο�_9��GX�����f�c�%�}�~�`�P���Y����l�N��Uʼ�
�!��&��)��������9��Q��A���%�n�u�u�>�����
����A��B��D���3�
�g�c�'�}�J�ԜY���F��h��6���
�!� �!�%��@ׁ�&����S��G_�����}�0�
�8�b�����I���F�_��U���0�_�u�u�w�}�;���&����l5��B�����b�
�e�3��o�N���B�����T������'�6� �2�l�B�������U��N�U���u�u�u�<��)�4���&����P��R1�@���3�
�g�a�'�}����Q����G��1����`�}�|�h�p�z�W������F�N��*����&�
�!�"�)����N˹��U��[����u�u�<�
�#���������F��V��A���
�a�e�%�w�`�}���Y���Z*��C1�����!� �!�'��j�(�������_��N�����&�9�!�%�n�;�(��M����O�I�\ʰ�&�u�u�u�w�}��������V9��E�� ���d�`�3�
�c�o���Y����9��h-�����'�6� �0�f�h�B���&����l��S��U���u�u�<�
�#���������F��V��M���
�g�a�%�w�5��������CP��Q��F���%�}�|�h�p�z�W������F�N��*����&�
�!�"�)����Aƹ��U��]����u�u�<�
�#���������F��V��M���
�g�a�%�w�`��������l��C�����0�}��6��<��������A�� _��E���
�g�l�%�~�p�����μ�e��h[�����a�b�|�n�w�}��������V9��E�� ���d�`�l�3��i�A���Y���F�N�����!��&�
�#�(����&����9��h]�@���u�=�;�}�2����&���� Q��G\��\��r�r�u�9�2�W�W���Y�ƥ�l��t��*��� �!�'�
�o��(���J����CU��N�����!��&�
�#�(����&����U��\�����h�_�u�u�w�}�;���&����l5��B�����b�
�e�3��o�N���Y����N��G1�*���f�c�
�g�g�}�W��PӃ��VFǻN��U����6�
�4�2���������S��h��F��
�f�_�u�w���������\��X�� ��c�
�g�i�w�)�(�������P�������1�<�
�<��/�;���&����T9��G��U���<�;�1�4��2��������]ǻN��9���1�
�0�8�f�m����K�֓�F���*���<�
�0�!�%�(�����θ�CW��Q��G���%�|�~� �$�:����&����l��1����b�|�n�u�w�4�(���¹��l4��P�����:�'�0�g�1��B���	���l�N��Uʴ�
�:�&�
�!�o�Gϩ�����V
��Z�*���f�b�
�g�g�}�W��PӃ��VFǻN��U���0�
�8�m�1��B���	��ƹF��{1�� ��� �
�e�
�"�n�N߁�K���@��[�����6�:�}�;�>�3�Ƿ�&����\��N� ���2�0�}��#�/�F���&����V9��S1�����
�
� �f�o��D���s���Z��1��*��
�g�i�u�f�}����Q����V��Z��Gӊ� �b�c�%�~�a�����έ�l��D��Ҋ�|�u�9�0�u��}���Y����9��hY�*��i�u�d�u�?�3�_�������^��^�� ��g�%�|�k�$�:����	����@��A_��E���0�&�u�e�l�}�WϷ�����]	��Q��A���%�u�h�}�4�-�(���K����CT��X�����;�!�9�d�f�f�W�������l ��Z�*��i�u�d�u�?�3�_���&����U��_�����u�%�6�;�#�1�E��Y����D��d��Uʼ�8�
� �a�g�-�W��[����[�������!�%�m�
�"�i�G���P����Z��SF��*���&�
�#�d�g�t����Y���9F���%���:�
�
��;���������l ��[�*��i�u�u�u�w�}��������lR��_��]���
�e�
� �d�m�(��I���W����ߊu�u�u�u��>�(�������F��E��Bۊ�g�3�
�a�n�-�L���Yӏ��T9��1��*���
�d�i�u��.����H���� U��G_�U���<�0�
�
�"�n�O���Y����l��^	�����f�
�d�_�w�}����&¹��lR��h�I���'�2��d�1��Bف�H����W	��C��F��u�u�9�
��(�O���	�����hX�����f�
�g�d�z�l��������l�N��*���d�m�
�d�k�}����O����U��h�D���d�1�"�!�w�t�}���Y����e9��Q��E���%�u�h�&�3�1��������AN��D�����%�6�;�!�;�h�(���Tӓ��Z��SF��'���9�
�
� �f�o�(��P���F��Y1��F���
�e�
�g�k�}��������E��X�����;�1�4�
�8�.�(���M���F��D�����
�0� �!�`�;�(��&���l�N�����c�3�
�d��n�K���Y���F��V ��*ي� �`�m�%�w�5����
����9��hZ�*��e�u�u�d�~�8����Y���F��h<�� ���b�3�
�e��l�}���Y����e9��h_�L���u�h�_�u�w�}�W���&����U��]�����=�;�}�&�2�����N���F�_��U���0�_�u�u�w�}�(�������l ��^�*��_�u�u�0��1�(���K����CU�
NךU���u�u�-�
�8�8����&����e9��h\�G���u�=�;�}�%�>��������
9��^��H��r�u�9�0�]�}�W���Y����V
��B1�Fފ�f�_�u�u�2��݁�����9��R�����u�u�u�-��2��������9��Q��@���%�u�=�;��0�(�������T��G��U��|�0�&�u�w�}�W�������\��C��*��
�
� �g�f��E�ԜY���F��@=��F���6�&�
� �e�l�(��E�ƿ�W9��P�����:�}�0�<�2�.����Q����V
��Q��C���%�|�g�|�l�W�W������� 9��h\�B���u�h�_�u�w�}�W���&����l��Z1�B���3�
�`�f�'�}����Q����G��1��*���`�%�}�|�j�z�P������F�N�����;�1�
�0�:�h�F�������T��UךU���0��9�
�"�o�@ځ�J���9F�N��U���
�:�0�!�%��Gف�&����V��G_�����}�8�
�g�%�:�C��Q���A��N�����u�u�u�u�1�-����&����lR��h8�� ��e�
�g�_�w�}����ƹ��lT��1��U��_�u�u�u�w�8�$���&����P��G]�����}�'�6�;��(�E��&���F�_��U���0�_�u�u�w�}��������V��Z��#���
�`�e�%�l�}�Wϰ�����l ��X�*��i�u�u�u�w�}��������l��C1��*��g�%�u�=�9�u��������lT��1��]���h�r�r�u�;�8�}���Y���U��Y��*���8�a�b��1��B���	��ƹF��R��ӊ� �g�e�
�d�a�W���Y�����V��Aۊ�0�
�e�b� �8�Wǭ�����R��B1�Gߊ�g�e�u�u�f�t����Y���F������d�
�0�
�n�o�}���Y����V
��B1�Fފ�f�i�u�u�w�}�Wϸ�	����V9��E��E܊�
� �g�e��l� ���Yە��l��^�����e�e�e�u�w�l�^ϻ�
��ƹF�N�����:�0�!�'��m�(�������9��d��Uʻ�"�<�;�<�����JŹ��Z�G1��؊�l�3�
�b�d�-�_������\F��UךU���0�&�2�7�#�o����K�ߓ� F������f�
� �g�f��E��Y����G	�G�U���;�"�<�;�>��(���K����CU�
N��#���
�d�3�
�o�j����Hӂ��]��_����u�0�&�2�5�)�C���&����l��S��*���g�`�
� �d�j�(��J�ƨ�D��]�N���u�;�!�6�%�$����K�ӓ�F�F�����;�<�
�
�"�o�Fց�JӉ��C9��D��*���;�!�3�
�e�d����s���\��X ��*���g�a�
�g�k�}��������l��hZ�Eʺ�u�6�%�
�2��G��B���	��T��G���
�`�f�%�w�`�_�������U��\�����'�:�
�:�3����M¹��]ǻN�����;�l�
�d�1��@ہ�K�����hX�����c�
�g�4�3�/�܁�����l��d��Uʺ�
�:�1�d�>�;�(��J����[�C��G݊� �d�d�
�e�<�Ϭ�¹��lW��1��\�ߊu�u�'�6�9�d�(�������9��R��]���
�a�3�
�a��EϿ�Ӕ��9��hV�*��n�u�u�:��2��������R��h�I���!�%�g�
�"�l�F؁�KӇ����h��D��
�g�n�u�w�2�(�������S��h�I���&�9�!�%�c�;�(��L����\��R�����
�0�
�e�`�f�W�������_	��1��*��b�%�u�h��/����&�ד�F9��X��Gʴ�1�!�%�b��(�F��&���9F������"�g�3�
�e�e����D�ή�^��R1��*���g�l�
�g�6�9����NŹ��lT��1��\�ߊu�u�#�'�;�*�D���&����l��S�����'�0�<�
�"�o�@ځ�KӇ����hW�����l�d�%�|�]�}�W�������lR��B1�Cߊ�g�i�u�7�:�/����&����S��G\�����8�
�b�3��l�G���P���F��R����� �d�`�
�e�a�WǼ�����l��B1�A܊�g�4�1�!�'�n�(���H����CT�=N��U���
� �d�e��n�K���Y���F��G1�����9�g�
���� ���Yۏ��V��R	��B��e�u�u�d�~�8����Y���F��G1�����9�g�
�n�w�}���&�ד�F9��]��G��u�6�'�,�f�;�(��O����R��e��ۊ�9�
�;�&�b�;�(��O����l�N��FҊ�g�3�
�d�e�-�W��Q����J9��Q��E���%�u�;�u�6�:�F�������@9��Q��D���%�|�_�u�w��O�������R��N�U¶�'�,�'�2�d�d�W���Y����Q��E��F��|�_�u�u�����Kʹ��Z�=N��U���u�%�6�;�#�1�Fׁ�?����D��F�����d�'�2�f�g�u�^��^���V
��d��U���u�4�
�:�$�����I���F��_��D���
�l�l�%�w�`�_����ԓ�_
��Y��F���
�l�d�%�w�3�W���&�ԓ�F9��Z��G��u�u�%�a��o����H�ޓ�F�F�����
�9�
�;�$�i����H�֓�F��SN����
� �f�g��o�L���YӖ��9��h��L���%�u�h�}�6�:�F�������\��h��L���%�u�'�'�!����K����l�N��Lߊ�
� �d�e��o�K���+����9��[1�����d�3�
�a�b�-�W�������F9�� _��G��u�u�%�l��l����I�Г�F�F����`�3�
�e�o�-�W���+����9��[1�����g�3�
�g��o�L���YӖ��9��Q��C���%�u�h�}�:��F݁�����9����'���0�
�9�
�2�2�(���H����CT�=N��U���m�<�
� �n�i����D�θ�C9��h��L���%�u�;�u�6�:�F�������\��h��L���%�|�_�u�w��O�������U��N�U¡�%�f�
� �f�j�(������R��1�����'�&�3�
�c�j����s���C9��D��*���;�!�3�
�e�d����D�θ�C9��1��*��d�%�u�:�w�-��������lW�=N��U���0� �!�g�1��Nׁ�K�����h8��*���`�a�%�u�9�}����Kǹ��lP��h�N���u�%��&�;��(���H����CW�
N�����2�6�#�6�8�u����ۓ��Z��SF�����
�e�g�%�~�h�^��Y����l4��B��B���
�e�
�d�k�}��������E��X�����0� �&�2�2�u����N����_��G]��@���n�u�u�%��.����&����^��G\��H���4�
�
� �f�n�(������^�� 1��*��`�%�|�_�w�}�(���K����^��Q��E���%�u�h�_�w�}�W���	����@��A_��D����"�0�u�5�0��������U��X�����|�h�r�r�w�1��ԜY���F��a��*���'�2�f�f�l�}�WϮ�/����P��B1�@܊�f�i�u�u�w�}�WϮ�/����9��O1��*��f�%�u�=�9�u��������U��[�����|�h�r�r�w�1��ԜY���F��[1�����3�
�e�f�'�f�W���	����9��h��D��
�f�i�u�w�}�W�������^��R	��M���"�0�u�&�;�)��������P��G��U��|�0�&�u�w�}�W���
����^��h��D��
�f�_�u�w�����H����U��h�I���u�u�u�u�6�����&����l^��^����u� �1�'�;�*�E���&����l��G��U��|�0�&�u�w�}�W���	����9��h��*��a�_�u�u��<�E��H����l ��^�*��i�u�u�u�w�}��������_��hY��3����"�0�u�5�0��������U��_�����|�h�r�r�w�1��ԜY���F��a��*���3�
�m�b�'�f�W���	����9��1�����
�g�g�%�w�`�}���Y���R��X ��*���g�b����}����Q����A��^1��*���f�l�
�g�g�}�W��PӃ��VFǻN��U���
�4�g�`��(�D��&����F�G1��؊�f�8�-�3��n�A���Y���F�N�����:�&�
�#�c�j�1���Y����N��Z�����<�
� �g�f��E��Y���O��[�����u�u�u�
�6�o�D߁�����R��N�����9�
�b�3��l�N���Y����K��R��*��
�
� �g�f��D�ԜY�Ƽ�e��h\�����d�l�%�u�j�.��������V��EF�����}�;�<�;�3�.��������V��EF�����}�
�4�g�e����Jʹ��F�D�����e�u�4�
�8�.�(���L����vO�N�\��u�u�%��;��N���&����l��S��*���g�g�
� �e�n�(��J�ƨ�D��_�N���u�%��9���O���&����l��S��U���u�u�4�
�8�.�(���K����V��N����� �1�'�9� �n����I�֓�N��S��D���0�&�u�u�w�}�WϮ�/����W��B1�L݊�g�_�u�u��<�E�������U��N�U���u�u�u�!�'�o�(���H����CW��_��]���
�
� �d�`��E��Y���O��[�����u�u�u�
��(�F��&����F�G1��؊�e�3�
�g�d�-�W��
����\��h����� �&�2�0������Kʹ��lT��1��\��� �&�2�0��0�(�������_��G����u�
�4�g�d�o�(���J����CU�
NךU���u�u�%�6�9�)���&����V�������;�0�3�:�����Aʹ��V�
N��R���9�0�_�u�w�}�W����ԓ� 9��h]�C���n�u�u�%��1�(܁�����9��R�����9�2�6�#�4�2�_���������V��G���
�d�f�%�~�v��������G��^�� ��g�
�d�|�]�}�W����ԓ�9��h\�E���u�h�_�u�w�}�W����ԓ� 9��O1��*��c�%�u�=�9�u��������9��C1��*��e�%�}�|�j�z�P������F�N�����9�
�
� �e�i�(��s���C9��[\��M���
�`�l�%�w�`�}���Y���]��R�����`�`�%�u�?�3�_�������l ��[�*��e�u�u�d�~�8����Y���F��O�����!�'�
�e�����Iʹ��l�N��#���
�
� �d�g��D��Y���F���*���3�
�d�l�'�}����Q����G�� 1��*��l�%�}�|�j�z�P������F�N�����!�%�`�3��o�A���B�����V��@ۊ� �g�l�
�e�a�W���&����P9��T��]���<�;�1�%��1�(�������Q��E�����;�1�!�%�n����@����O��N�����9�
�f�3��m�A���Y����G��X	��*���!�'� �&�0�8�_����ԓ�9��P1�G���~� �&�2�2�u����M���� V��h�\�ߊu�u�
�4�e�h�(���J����CU�
NךU���u�u�
�4�e�o�B������� T��h����u� �1�'�;�*�C������� T��h�E���u�d�|�0�$�}�W���Y����l0��1��Gڊ� �f�g�
�d�W�W���&����lS��1��*���e�%�u�h�]�}�W���Y����V
��Q��@���%�u�=�;��/����K����S��h�E���u�d�|�0�$�}�W���Y����V��[Z�� ��b�
�f�_�w�}�(���K�ӓ�F9��^��F��u�u�u�u�w�<�(���
����R�������8�
�
�0��j�E��Y���O��[�����u�u�u�%�4�3����Kǹ��V��d��Uʥ��9�
�
�"����I����Z�=N��U���u�%�6�;�#�1�Eہ�?������YN�����2�
�
�
�"�l�@ց�K���F�G�����_�u�u�u�w�����M����lU��UךU���
�4�g�c�1��A���	�����h�����0�!�'� �$�:����&����l_��B1�F܊�f�u�u�;�>�3�Ǫ�	����U��X�����n�u�u�%��1�(؁�����9��R�����u�u�u�-��2��������9��Q��@���%�u�=�;��/����&����T��G\��\��r�r�u�9�2�W�W���Y�Ƣ�D5��h��G��
�f�_�u�w�����A����P��h�I���u�u�u�u�9�*��������U��N�����:�
�:�1��(�E��&���F�_��U���0�_�u�u�w�}��������lT��1��N���u�%��9�����JŹ��Z�=N��U���u�8�
�d��8�(��Iӑ��]F��Z��G���2�f�g�}�~�`�P���Y����l�N��Uʥ�f�3�
�c�n�-�L���YӖ��R
��D1�*���f�a�
�f�k�}�W���Y����l0��1�D���-�3�
�e�d�-�W����ι�W��[��F���!�3�
�e�`�-�_���D����F��D��U���u�u�%��;��(�������W��UךU���
�4�g�&�1��G���	���l�N��Uʴ�
�:�&�
�!�e�Gϩ�����^��1����d�}�|�h�p�z�W������F�N��*���&�
�#�m�e�m�G�ԜY�Ƽ�Z*��C1�����:�
�4�!�1��B���	�����h�����0�!�'�'�$�'�_���������{1��*���
�:�%�&�1��B���	���O�=N��U����9�
�:��2��������Q��N�U���u�u�u�4��2�����ד���YN�����c�
� �f�f��D��Y���O��[�����u�u�u�8��k�(���J����CW��N�����!�<�
� �e�k�(��E����V
��R
�����
�
� �g�d��DϦ�Ӈ��P	��C1��D��n�u�u�%�9�)�݁�����9��R��]���0�0�
�0�8��(���J����CU��X�����;�!�9�d�f�f�W���	����l��B1�MҊ�g�i�u�1�;�)��������l��hZ�Gʭ�'�4�
�:�$��ށ�P���F��X�����c�
�g�i�w�)�(�������P�������1�!�%�d�g�;�(��&���F��D�����%�6�;�!�;�k�F���s���C9��h��A���%�u�h�&�3�1��������AN��D�����8�
�a�3��m�(��Y�ƹ�@��R
�����;�!�9�c�f�t�}���Y����U��_�����h�_�u�u�w�}��������EU�������8�
�g�'�0�i�E���P���A�R��U���u�u�u�4��2��������9F�N��U���d�d�6�&��(�@���	�����h�����0�!�'�'�$�'�_�������\��1��*��
�g�y�g�~�W�W���	����9��hY�*��i�u�!�
�8�4�(�������]��Y��3؊�
� �`�m�'�t�\ϫ�
����WN��h�����#�g�g�|�]�}�W���Y����l��C1��*��c�%�u�h�$�9��������G	��E�����<�;�1�%�$����J¹��J��G����u�:�d�3��n�F���Y����G��X	��*���!�'� �&�0�8�_�������^��E�����;�1�4�
�8�.�(���K���l�N��Uʥ�&�
�
�4�#�;�(��&���F��S1�����#�6�:�}�2�4�ǭ�����C	��h_�� ��m�%�|�f�~�f�}���Y����lW��B1�M���u�h�&�1�;�:��������F��P ��]���d�3�
�g��o�W�������V��G1�����9�d�
�|�l�}�W���YӖ��9��D�� ��a�
�d�i�w�)�(�������P�������&�2�0�}�8�o����J�֓�O�G����u�%�&�
�"�l�C߁�K���@��[�����6�:�}�;�>�3�ǘ�&���� Q��N�� ���2�0�}�%�4�3����H����]ǻN�����3�
�f�
�d�a�W���Y�����R	��*���a�a�%�u�?�3�_���&�֓�F9��1��]���h�r�r�u�;�8�}���Y���G��_�����f�
�f�_�w�}����
����9��h_�B���u�h�}�
�����H¹���������d�a�%�|�]�}�W�������]9��Q��C���%�u�h�}���F���&����l��V �����
�0�
�m�g�f�W�������@��h[�� ��e�
�g�i�w�/����&����_��G\�����7�!�3�
�f�n����s���B��D�����3�
�m�m�'�}�J���&����l ��V�*��4�1�$�<������I���9F������2�
�
� �d�k�(��E����l��1��*��g�%�u�;�w�?��������T��d��Uʤ�
� �d�`��n�K���Y���F��D ��*���
�b�b�"�2�}����H����lW��1��]���h�r�r�u�;�8�}���Y���G��V�� ��a�
�f�_�w�}��������U��N�U���4�g�g�
�"�o�Dց�K����\��XN�N���u�'�d�3��l�(��E����^��1��*��
�g�4�1�#�-�Bف�����l��d��Uʧ�g�3�
�d�b�-�W��[����[����*��
� �g�b��l�JϿ�&����G9��1�U���0�w�w�_�w�}�(܁�����9��R��W���"�0�u�!�'�l�@�������F�V�����
�#�d�e�w�1����[���F��1��*��b�%�u�h�u�� ���Yے��lW��h��*��a�h�4�
�8�.�(���H���V
��L�N���u�'��d�1��N߁�K���@��[�����6�:�}�=�1�����Q����T�������!�9�`�
���1���?����J��h�����}�;�<�;�3�z�P�������9��hV�*��f�x�u�:�9�2�G���P��ƹF��h8��*���g�b�
�g�k�}��������E��X�����1�!�%�m��(�E��&���F��P ��]���
�a�3�
�a�i����B�����h[�� ��l�
�g�i�w�)�(�������P�������!�%�m�
�"�o�Oہ�H���@��R
�����c�3�
�c�o�-�^��Y����l0��B1�Fӊ�g�i�u�!��2����������Q�����}�;�<�;�3�<�(���
����R��q(��3������y�8�4����ۓ��Z��SF��R��!�%�g�
�"�l�Eց�H����F��@ ��U���|�|�_�u�w����@����Z���*���3�
�d�d�'�}��������l ��_�*��n�u�u�'�>�4�(���H����CT�
N�����g�
� �d�b��Fϱ�Y����A��V�\�ߊu�u�
�
�e�;�(��N����[�C��D���3�
�d�l�'�}�Ϭ�K����W��h�N���u�'�<�<��(�E��&���F��Z��Aӊ�0�
�e�b�8�}�(܁�����9��UךU���
�
�a�3��m�E���Y���G��[�����a�a�u�'�%�i����I�ѓ�O��N�����<�3�
�g�f�-�W��Q����P��B1�E݊�d�:�u�
�"�l�N܁�K��ƹF��R�����a�d�%�u�j�u����Iʹ��lW��1��U���u�%�6�;�#�1�F��B�����1��*��
�g�i�u�#�-�F�������9����U���6�;�!�9�f�l�L���YӔ�� 9��hV�*��i�u�!�%�f�i����Lǹ���������!�9�d�d�l�}�WϬ�Ĺ��lT��1��U��}�:�9�-����������l)��r�����3�
�f�m�'�}����	����@��A_��\�ߊu�u�0�m�1��C���	���N��G1�L���2�a�c�u�8�}��������EW��UךU���0�l�3�
�b�n����D�θ�C9��1��*���`�%�u�:�w�-��������lW�=N��U���
� �d�b��o�K�������P��B1�Cي�f�-�'�4��2����¹��l�N�����%�e�3�
�b�j����D�θ�C9��1����c�u�;�u�2�d����L�Փ�O��N�����!�%�d�3��o�G���Y���@��C��*���d�`�
�g�6�9����O����lW��1��\�ߊu�u�0�
�:�l�C�������Q��h�I���&�9�!�%�e�;�(��K����K	��V�����
�#�
�|�]�}�W���&����9��h_�C���u�h�_�u�w�}�W����ԓ�l ��\�*��"�0�u�&�;�)��������V��F�U���d�|�0�&�w�}�W���Yӕ��l��1��*��d�%�n�u�w�.����	�Փ�F9�� Z��G��u�!�%�c��(�F��&����\��G1�����9�d�d�n�w�}��������l ��\�*��i�u�&�9�#�-�(���H����CT��Y
�����8�d�
� �f�j�(��B�����h��Dߊ� �d�m�
�d�a�W���Y�����V��F���
�g�b�%�w�5��������CW��Q��G���%�}�|�h�p�z�W������F�N�����%�g�3�
�e�k���Y����V
��Z�F���8�'�4�
�"�o�N܁�K�����h]�����f�d�u�'�>�0�E�������O��N�����!�%�c�3��o�C���Y���D��_��]���;�1��
�2��@��Y�ƿ�T�������!�9�d�
�a�t����Y���9F���*���d�l�1�8�%�<�(���K����CT�
N�����
� �g�g��o�����ѓ�F9��V��G��u�u�&�9�#�-�@���&����l��S�����!�%�c�3��o�C���Y����G��1��*��g�%�|�_�w�}��������l��X�����
�a�m�%�w�`�_���&����_��R�����3�
�a�a�'�}�Ϫ�	����U��]�����_�u�u�0��0�Fׁ����� 9��R��]���
�e�
� �f�k�(���Ƹ�C9��h ��*���d�e�
�g�l�}�Wϭ�����_��B1�Dӊ�g�i�u�!�'�n�(���H����CT��Y
�����8�d�
� �f�l�(��B�����h��D���
�g�l�%�w�`�_���&¹��lW�� 1��U���u�%�6�;�#�1�F��B�����h��Gڊ� �d�g�
�d�a�W���Y���4��P�����:�0�
�
�"�l�N؁�Kӑ��]F��R����
� �d�d��o�G���Y�����RNךU���u�u�0�
�"�l�@ށ�K���F��[1�����3�
�`�d�'�}�J�ԜY���F��Y	��*���
�0�:�
�"�l�@؁�Kӑ��]F��R����
� �d�d��o�G���Y�����RNךU���u�u�
�`�>�;�(��H����9F���*���g�
� �d�g��E��Yے��lT��E��F��u�:�u�%�4�3����H���9F���*���g�
� �d�f��E��Yے��9��h_�A���u�;�u�&�2�����N���9F���*���g�
� �d�e��E��Yے��lT��E��F��u�;�u�&�2�����N���9F���*���g�
� �g�e��D��Y���F������`�3�
�e�g�-�W����θ�C9��h��G��
�g�e�u�w�l�^ϻ�
��ƹF�N��*���g�a�'�2�d�m�L���Yӕ��l��X�����'�4�
� �d�n�(��E����^��1��*��l�%�u�'�#�-�F�������R��G�U���&�9�!�%�a�;�(��J����[�N��U���&�9�!�%�b�;�(��K����D��F�����%�b�1�8�%�<�(���K����CT�N��R��u�9�0�_�w�}�W���&����lR��R	��L��_�u�u�0��0�E�������T��Q��F���%�u�h�}�2����N����\��Y1��*��m�%�u�'�#�-�F�������_��G�U���&�9�!�%�`�;�(��I����[�C��C���2�f�b�u�8�}��������EW��UךU���0�
�8�g��(�E��&���F��Z�����e�`�%�u�9�}��������V��d��Uʦ�9�!�%�l�1��Fف�J���9F�N��U���
�d�
� �b�m�������G��_�� ���a�%�}�|�j�z�P������F�N�����:�&�
�#�o�m�}���Y����G��h��F��
�g�i�u�f�}����Q����Z9��E1�����
�0�
�e�w�}��������ET��N�����e�n�u�u�$�1����I����T��G\��H���8�
�d�3��k�(������C9��Y�����d�n�u�u�$�1����H����U��G\��H��� ����f�;�(��&����]��R����
� �b�a�'�t�}���Y����G��1��*��g�%�u�h��8�(���J¹��T9��[�����8�
�g�
�"�l�C݁�J��ƹF��R����
� �d�m��n�K���Y���F��h8��G���3�
�c�m�'�}����Q����G��1��*��g�%�}�|�j�z�P������F�N�����!�%�l�'�0�n�B��Y����V
��Z�*���d�l�
�g�k�}����H�Г�F9��\��Fʭ�'�4�
�:�$��ށ�P���F��[1�����3�
�b�e�'�}�J�������CU��E��F���u�;�u�0��0�Dہ�����9��UךU���0�
�8�f��(�F��&���FǻN��U���
�4�g�c�1��A���	�ƻ�V�D�����`�3�
�b�g�-�_���D����F��D��U���u�u�&�9�#�-�D���&����l��=N��U���
�8�f�
�"�j�E���Y���Z��1��*��
�g�4�1�#�-�Cہ�����l��d��Uʦ�9�!�%�m�1��Aہ�K�����h_�*���m�a�%�u�%�)���&����U��V��G��u�u�&�9�#�-�N���&����CT�
N�����m�3�
�a��o����
����^��h��L���%�|�_�u�w�8�(���J����T��h�I���u�u�u�u�#�-�Fց�����9�������8�
�
� �f�k�(��I���W����ߊu�u�u�u�'�>��������]ǻN�����8�a�
� �n�k����D���F�N�����
�9�
�;�$�n����M˹����YN�����8�f�
� �n�m����P���A�R��U���u�u�u�'�!����K����9F���*���a�
� �l�e�-�W��s���F�e��ۊ�9�
�0�:�����A����D��F�����%�l�3�
�`��E��Y���O��[�����u�u�u�
�b�4�(���@�ԓ�]ǻN�����8�a�
� �f�m�(��E����^��1����b�u�:�u�'�>�����ד�]ǻN�����8�a�
� �f�l�(��E����^��h��D��
�g�4�1�>�3��������V��d��Uʦ�9�!�%�a�1��O���	���N��G1�*���
�m�a�4�3�4����H����lU��G�U���&�9�!�%�b�;�(��O����[�N��U���%��9�
��(�E��&����[����*���3�
�e�g�'�u�^��^���V
��d��U���u�%��9��d����J����9F���*���a�
� �g�n��D��Y���F���*���a�
� �g�o��Dϩ�����V
��Z�F���8�'�4�
�"�o�N܁�K���F�G�����_�u�u�u�w�����Hʹ��T9��W�U���&�9�!�%�`�;�(��M����[�C��FҊ�0�
�m�b�/�/��������_��G�U���&�9�!�%�o�;�(��M����[�C��G���
�d�l�%�w�3�W���	����T9��V����u�0�
�8�c����L����Z���ي� �g�g�
�e�%�Ͽ�&����G9��1�N���u�&�9�!�'����MŹ��Z���*��
� �f�e��o��������A��_�\�ߊu�u�0�
�:�h�(���K����CT�
N�����3�
�a�m�'�}��������CR��Q��A���%�|�_�u�w�8�(���L¹��lT��1��U��}�:�9�-����������l)��r�����3�
�f�m�'�}��������l��h��G��
�g�n�u�w�.����	�ԓ�F9��\��G��u�!�%�b��(�E��&����]��R�����
� �g�b��o�L���Yӕ��l��]�� ��l�
�g�i�w�.����	����W��E	��*���g�m�
�g�/�/��������_��G�U���&�9�!�%�c�;�(��L����[�C��Mڊ�0�
�e�m�6�9��������l��hZ�G��u�u�&�9�#�-�B���&����l��S��U���u�u�4�
�8�.�(���&�ƻ�V�D�����e�'�2�a�d�u�^��^���V
��d��U���u�4�
�:�$��܁�B�����h��@܊� �g�a�
�d�a�W���Y�����h��@ߊ� �g�f�
�d�*��������]��Q��@���%�}�|�h�p�z�W������F�N�����
�`�m�%�l�}�Wϭ�����Q��B1�@ފ�f�i�u�u�w�}�WϿ�&����G9��1����u�&�9�!�'�i����L�ӓ�N��S��D���0�&�u�u�w�}�WϿ�&����G9��1����u�0�
�8�b����H˹��Z���*���3�
�g�l�'�}����	����@��A_��\�ߊu�u�0�
�:�h�(���&����P��G\��H���0�
�8�d��(�F��&����\��G1�����9�d�d�n�w�}��������l ��]�*��i�u�!�%�f�m����K�ғ�F��SN�����%�m�3�
�d�e����s���@��C��*���f�`�
�f�k�}�W���Y����l��[�����:�%�6�&��(�D��&����[����*���a�3�
�`�a�-�_���D����F��D��U���u�u�<�
�2�4��������l ��h"�����3�
�`�l�'�f�W���
����^��h��F��
�g�i�u�$�1����OĹ��^	��V �� ��f�
�g�-�%�<�(���
����9��d��Uʦ�9�!�%�d�1��D���	���N��G1�D���
�g�l�%�w�3�W���&����9��h]�A���|�_�u�u�2����&���� Q��G\��H���0�
�8�g�c�9��������lU��1��U���u�%�6�;�#�1�F��B�����h��Cي� �f�b�
�e�a�WǪ�	����l ��\�*��4�1�&�9�#�-�E���&����l��d��Uʦ�9�!�%�
�"�n�Bց�K�����h_�*���f�e�
�g�/�/��������_��G�U���&�9�!�%��(�D��&���F��R�����a�l�u�;�w�8�(���O���� S��h�N���u�&�9�!�'����Nù��Z�=N��U���u�;��'�8��W����ο�_9��GY�� ��c�
�g�e�w�}�F�������9F�N��U���
�8�`�3��h�F���B�����h��L݊�0�:�2�;�1��G���	���N��G1�����f�b�u�'�>�0�(���&����]ǻN�����8�l�3�
�e�h����D�Ν�r(��y-�����b�g�4�1�$�1����&����R��G\����u�0�
�8��(�D��&���F�N�����<�
�<��%�����&���� V��
N��*���&�
�#�
�~�8����I��ƹF�N�����!�d�6�&��(�B���	�����h�����0�!�'�'�$�'�_�������[9��C1�����`�
�f�y�e�t�}���Yӕ��R��1��*���
�f�i�u�w�}�W�������
9��h[�*��"�0�u����9���&���� R��F�U���d�|�0�&�w�}�W���YӒ��lR��Q��A܊�g�_�u�u�w�}��������G9��h_�F���u�h�&�1�;�:��������A��M�����1�&�
�8��(�F��&��� T�dךU���=�4�!�3��m�A���Y���F�N�����l�3�
�e�a�-�W����Ν�r(��y-�����b�g�e�u�w�l�^ϻ�
��ƹF�N�����
� �d�`��o�}���Y����l��^	��D���
�m�b�%�w�`�}���Y���G��W�� ��l�
�g�"�2�}��������l ��V�*��e�u�u�d�~�8����Y���F��R����
� �d�d��o�}���Y����l��^	��D���!�3�
�m�f�-�W��Q����l��^	��D���
�m�b�%�w�2�W�������l
��h_����u�<�;�4�$�:�(���H����CU�
NךU���u�u�8�
�d�;�(��@����D��F�����%�a�3�
�n�i����P���A�R��U���u�u�u�&�;�)��������_��UךU���<�;�4�&�0���������9��R��]���;�4�&�2��(�F��&����\��G1�����9�d�d�n�w�}��������F9��[��F��u�
�4�g�e����Jʹ��U��S�����a�n�u�u�#�-�G���&����l��S�����<�;�<�
��(�F��&����]��R����
� �d�e��o�L���YӒ��W��B1�M݊�g�i�u�:�2�;����&����S��G\��ʦ�2�
�&�<�9�l��������W��G�U���!�%�g�3��l�N���Y���Q��E	��*���
�l�b�4�3�.����	�ѓ�F9��Z��G��u�u�!�%�d�;�(��L����[�Y�����<�
�
�0��d�Gϱ�Y����P��B1�Bӊ�g�n�u�u�#�-�C���&����l��S�����g�
�0�:�0�3����@�ޓ�F��EN��*���&�
�#�
�~�W�W�������U��\�����h�}�'�0�0�i�(�������l��Q��L���%�u�'�!�'�d�(���K����CT�=N��U���d�
� �f�o��E��Yے�� T��S�����
� �f�b��o��������]��[��D��u�u�!�%�`�;�(��I����[�U�����e�1�8�'�6��E���&����l��X�����b�3�
�d�g�-�^�ԜY�Ƹ�CW��Q��G���%�u�h�&�3�1��������AN��D�����
�4�g�`��8�(��N���F��P ��]����'�:�
�~�f�W�������U��_�����h�}�8�f�n�9��������lW��1��U���u�%�6�;�#�1�F��B�����1��*��d�%�u�h������J�ѓ�F��SN�����
�f�d�%�~�W�W�������l��X�����
�f�f�%�w�`�_���&�ԓ�F9��]��Fʺ�u�0�
�8�f����@ʹ��]ǻN����e�6�&�
�6�)����KŹ��Z�=N��U���u�%�6�;�#�1�F݁�Y����N��v ��;��� �f�e�%��t�J���^�Ʃ�@�N��U���4�
�:�&��+�E��s���G��X�����2�;�3�
�`�d����D�θ�C9��1��*��a�%�u�'�$�1����N����lU��G�U���!�%�d�
�6�)����&����^��N�U���u�u�u�4��2�����ԓ���YN�� �����d�3��n�(��I���W����ߊu�u�u�u�'�>��������]ǻN����f�1�8�'�6����I˹��Z���M���3�
�g�a�'�}�ϼ�����V��R�����<�3�
�f�c�-�^�ԜY�Ƹ�CU��h
�����;�3�
�l�o�-�W��Q����l��Q��L���%�u�'�7�:�/��������T��^_�� ��l�
�g�n�w�}����KĹ��^	��V �� ��b�
�g�i�w�-�Dׁ�K���� W��h����'�0�2�a��8��������U��Y�����_�u�u�8�d�;�(��H����[�D�����b�3�
�g�n�-�W���
����^��h ��*���d�c�
�g�l�}�WϪ�	ǹ��lW��1��U��}�0�&�2�5�)����J����R��D�����g�3�
�l�c�-�^�ԜY�Ƹ�CS��B1�Lۊ�g�i�u�:�2�;��������9�������
�&�<�;�9�)����@�ӓ�O��N�����
� �g�a��o�K�������T��B1�L݊�g�4�1�&�;�)��������V��G�U���!�%�
� �f�o�(��E����^��1�����4�
� �d�f��EϦ�Ӈ��P	��C1��D��n�u�u�!�'����K����[�[*��*���m�m�%�u�9�}��������9��UךU���8�l�3�
�`�k����D�ο�_9��G]�����f�c�u�'�$�1����Kǹ��G9��h_�E���|�_�u�u�:��G߁�����9��R��W���"�0�u� ��.�4���&����P��R1�M���2�a�c�u�w�-��������lT�R��U��n�u�u�!�'�l�F���&����l��S��D���=�;�}��4�����*����G��h_�*���
�e�f�h�6�����&����O��[��W���_�u�u�8��m�(���J����CT�
N��Wʢ�0�u� �
�$���������F��Z�����a�c�u�u�'�>�����Փ�F��D��E��u�u�!�%�f�n����L�֓�F�L�U���;�}�<�;�3�4�(���:����`��T����d�d�
� �d�e�(��Y�ƿ�T����%���:�
�|�u�;�8�U���s���G��^�����`�`�%�u�j�4�(���;����lT��h��F��
�g�f�u�8�3���B�����h_�*���d�c�
�f�k�}�������� W��F�U���;�:�d�|�]�}�W���&����U��^�����h�%�&�
�"�l�C߁�K����W	��C��D��u�u�u�u�#�-�F߁�����
9��R�����9�2�6�#�4�2�_�������Z��SF����
� �d�b��l�[��P��ƹF��Z��D؊� �d�e�
�d�a�W���H����U��h�D���:�;�:�d�~�W�W������� 9��hZ�*��i�u�'�2��l����LŹ��P��N����!�u�|�_�w�}����Hƹ��lR��h�I���'�2��d�1��Bف�H����F��S�����|�_�u�u�:��Fف�����l��S�����
�
� �`�c�-�_��T����\��XN�N���u�!�%�d�`�;�(��&���F��G1�*���`�e�%�}�o�p�FϺ�����O��N�����d�m�3�
�f��F��Y����_��B1�A���}�m�x�d�3�*����P���F��G1�L���
�f�
�f�k�}����&Ź��lS��h����;�0�0�}�9�4��������9��D�� ��c�%�|�u�8�3�Ϫ�&����T��B �����}�8�
�c�4�.�(���O�Г�O������:�<�!�2�%�(�����θ�C9��h�����
�g�
�d�~�`�GϿ�Ӓ��Z��P�� ���2�0�}�8��k����&����P��G�H��u�9�0�w�u�W�W�������l ��_�*��i�u�!�
�8�4�(�������[��h�� �&�2�0�}�:��G���&����l�������2�'� �&�0�8�_��Y�ƿ�l��h�����
�e�f�%��l�FϺ�����O�G�U���!�%�d�e�1��Aہ�H���G��Z�� ��g�%�}�u�w�}�������9F���*��
� �c�a�'�}�J�ԜY���F��h�����#�
�c�"�2�}����Lƹ��lP��h�E���u�d�|�0�$�}�W���Y����l	��h��C���%�n�u�u�#�-�F�������9��R�����9�2�6�#�4�2�_�������]��Y�����d�d�3�
�`��D��M����F�C��D���3�
�m�
�e�a�W���&����P9��T��]���3�
�0�!�"�.����Q����\��h��A���������^ê�&����T��B �����}�e�u�u�:��E݁�����l��_��U���;�:�e�|�~�f�W�������R��B1�G���u�h�}�8��o�(���O�Г�F��EN��*���&�
�#�a�d��1���?����uO��N�����d�c�3�
�a�o����DӖ��R
��1��*��c�%�}�b�3�*����N��ƹF��Z��G݊� �d�`�
�f�a�W����ԓ�l ��X�*��d�x�d�1� �)�W���s���G��\�����c�a�%�u�j�-�!���&Ź��lW��1��]��1�"�!�u�`�f�W�������_��B1�C���u�h��
��(�B���	������Y��A��u�u�!�%�f����J¹��Z�_�����u�&�2�0��0�(ց�����9��N����0�}�%�6�9�)���&�����RN��W�ߊu�u�8�
�d����K����[��Z��L���
�c�
�g�f�}�������9F���*��
� �m�a�'�}�JϮ�
¹��U��V��G��u�:�;�:�f�t�}���Y����U��Q��@ފ�f�i�u�:�e�l����@˹��W��S�����d�n�u�u�#�-�F�������^��N�U���d�d�3�
�o��E��Y����G	�G�U���!�%�d�l�1��F���	�����V��G݊� �g�f�
�e�d�Z������\F��d��Uʡ�%�d�
� �d�i����Dӏ��T9��Q��FҊ�d�`�u�u�w�2����I��ƹF��Z��Aڊ� �g�m�
�d�a�W����ԓ�9��h\�L���}�f�1�"�#�}�D��Y����^��_�� ��m�
�f�i�w�����KĹ��lT��1��]��1�"�!�u�g�f�W�������U��B1�@Ҋ�f�i�u�
�6�o�Cށ�����9��\����!�u�f�n�w�}����H�ғ�F9��Z��F��u�7�:�
��$��������A9��h+�����
� �g�l��o�Qϼ�����vV��C1�����'��
�$�6��(���K����CT�=N��U���
�a�
� �e�i�(��E�ƪ�C9��b"��:����9�<�9��o�(�������9��\�X��1�"�!�u�~�W�W�������l ��_�*��i�u�!�
�8�4�(�������]��Y��3؊�0�
�b�e�w�}��������C9��Y����
��|�n�w�}����H�ғ�F9��\��D��u�-�
���$��������_��Y��*���g�d�
�g�e�}�W�������V�=N��U���
�`�3�
�f�l����D������YN�����1��
�0��j�G���Y����V��G1�����9�d�
�b�~�8����I��ƹF��Z��Cڊ� �f�l�
�f�a�W�������@��C�����
�b�
�g�1��C���	����K�
�����e�n�u�u�#�-�F�������S��N�U���6�
�4�0��/��������lW��Q��A���%�}�d�1� �)�W��B�����h_�*���f�d�
�f�k�}�;���&����l5��B�����b�
�g�3��i�N���Q����\��XN�\�ߊu�u�8�
�a�;�(��&���F��S1�����#�6�:�}�9�4����?����lU��h�U���;�<�;�1�6�����&����l ��G�U���!�%�d�
�"�i�E���Y���D��_��]���;�1�!�%�f����O����X��^	��´�
�:�&�
�!�o�D���Y����D��d��U���u�!�%�d��<����&����l��S�����:�<�
�0�#�/�����ο�T����*���3�
�d�b�'�t�D���B���F��G1�*���d�m�
�g�k�}�G������C9��D��*��� �d�m�
�e�`��������_��h^�����u�d�n�u�w�)���&����Q��G_��Hʸ�;��3�
�g�d����M�����Y��E��u�u�!�%�f�;�(��N����[�L�����}�g�'�2�d�e�W���	����@��A_��D���0�&�u�e�l�}�WϪ�	����U��\�����h�&�1�9�0�>�����ξ�@�������1�$�
�&�>�3�F���&����l��\�\�ߊu�u�8�
�f�;�(��&���F��S1�����#�6�:�}�9�4��������9��D�����3�
�g�
�d�}�W���������h8�� ��m�%�|�n�w�}����K����lW�� 1��U��w�w�"�0�w�.����Q����l ��]�*��u�u�<�;�3�<�(���
����T��G�����u�e�n�u�w�)���&����_��G_��Hʡ�%�m�3�
�g�o����M�����Y��E��u�u�!�%�e����NĹ��Z�D�����6�#�6�:��8��������]��G��*���!�3�
�f�a�-�^��P��ƹF��Z��@���
�d�l�%�w�`����H¹��lW��1��]��x�d�1�"�#�}�^�ԜY�Ƹ�C9��h��D��
�g�i�u�#�����&����\��_��*���=�}�<�;�3�0�������� _��G�����!�2�'� �$�:����I���G��Z�� ��b�
�d�f�z�}�������O�=N��U���
�b�3�
�c�j����D������YN�����1�%�&�
�"�l�C߁�K���@��R
�����;�!�9�d��k�^ϻ�
���]ǻN�����m�3�
�d�a�-�W������l ��^�*��!�
�;�0�2�u��������^��1����� �d�a�
�f�t�����Ƹ�l��R	��]���<�;�1�!�'�l�(�������W��h�\���=�;�}�:�>�)��������]��C��DҊ�4�!�3�
�f�o����G����R��C�����0�}�;�<�9�9����H˹��@��B1�A؊�d�|�h�f�w�1����[���F��G1�*���d�g�
�d�k�}��������E��X�����0� �&�2�2�u��������U��Z�����`�|�n�u�w�)���&����U��^�����h�}�8�
�`�;�(��N����K	��V�����
�#�
�|�]�}�W���&����lU��h�I���!�
�:�<��8��������VN��D�����-�
�8�
��(�D���	���O�=N��U���
�e�3�
�c�l����D������YN�����g��d�3��i�D���Y�ƭ�l��D�����e�u�9�0�u��}���Y���� W��B1�Mӊ�g�i�u�d�w�5�����ԓ�F9��^��G��4�
�:�&��+�E��PӃ��VF�UךU���8�
�g�3��m�@���Y���G��1����b�u�'� �3�/��������U��G�U���!�%�f�
�"�l�Nց�K���4��P�����:�0�
�
��i����J����K	��V�����
�#�
�|�]�}�W���&�ғ�F9��1��U��!�%�d�
�"�n�A���Q���F��@ ��U���_�u�u�8��h����@�ד�F�F�����'�2�f�`�w�2�W�������l
��h_����u�8�
�c�1��O݁�H���@��[�����6�:�}�0�>�8��������V��C��#���3�
�b�
�c�q�E���s���G��Y�� ��c�%�u�h��-��������lW���*��
� �a�g�'�t�}���Y���� ^��B1�G���u�h�w�w� �8�WǪ�	����l ��X�����u�%�6�;�#�1�A܁�PӃ��VF�UךU���8�
�l�3��i�(��E�ƿ�W9��P�����:�}�;�<�9�9�1݁�&����^��G��U���<�;�1�4��2�����ԓ�uV�d��Uʡ�%�f�3�
�c��F��Y����l0��B1�M���}�f�x�d�3�*����P���F��G1�*���`�c�%�u�j�.��������V��EF�����0�}�%�6�9�)���&���F��D�����g�d�3�
�e��E���s���G��_�� ���a�%�u�h�u�� ���Y۠��9��h[�*��h�4�
�:�$�����H����_��^�����u�8�
�g�1��@ہ�K���W�@��U �&�2�0�}�?�<��������9��N� ���2�0�}�%�4�3����H����O��[��W���_�u�u�8��n����H˹��Z�=N��U���u�%�6�;�#�1�A��Y����N��G1�*���a�g�%�}�~�`�P���Y����l�N��Uʥ�:�
� �a�e�-�L���YӒ��lR��Q��Mڊ�g�i�u�d�w�5��������V��_1�����3�
�`�
�d�}�W���������T�����d�
�g�|�2�.�W��B�����hZ�����m�
�d�i�w�)�(�������P������� �&�2�0��5����H����G9��h[�*��y�a�|�_�w�}����O����_��G\��Hʦ�1�9�2�6�!�>��������A��CF�����}�4�
�
��(�B���	����\9��C�� �&�2�0�}�g�}�W���&�ӓ�F9��1��]��d�1�"�!�w�t�^���s���F�C��A݊� �c�e�%�w�`��������l��C�����/�}�<�;�3�)���O����Q��G_��F���n�_�u�u�:��O���&����l��S�����:�<�
�0�#�/�����ι�@��R
�����f�'�2�f�n�t�B���B�����hZ�����e�
�g�i�w�)�(�������P�������0�!� �&�0�8�_���&�ѓ�F9��1��\ơ�
�;�0�0��3��������@��_1�����6�&�
� �b�m����H����\��XN�\���n�u�u�!�'�i����I�Г�F�L�U���;�}�;�<�9�9��������lW��1��\�� �&�2�0��-��������9��G�����w�w�_�u�w�0�(�������9��R��W���"�0�u�&�0�8�_���&�ߓ�F9��1��\��&�2�0�}�'�>�������� P������w�_�u�u�:��F���&����l��S�����:�<�
�0�#�/��������GN��D�����%�6�;�!�;�h�(ܘ�?����u ��q(�����;�0�0�}�9�4����^�����hZ�����d�c�%�}�f�l��������O�d��Uʡ�%�`�
� �a�m����Dӕ��l
��^�����'� �&�2�2�u�E�������9��N�� ���2�0�}�%�4�3����H����uO�=N��U���
�f�3�
�c��E��Y���D��F�����}�g�d�3��o�(��Y�ƿ�T�������!�9�d�
�f�t����Y���9F���*���3�
�`�
�e�a�W���&����P9��T��]���<�;�1������A����M��Y�����4�
�:�&��+�E���<����F�C��@ߊ� �c�m�%�w�`�U���������Y�����`�
� �c�e�-�^���
����WN��h�����#�g�f�|�w�1����[���F��G1�*���b�a�%�u�j��Uϩ�����l4��B��G���
�l�
�g�j�<�(���
����R��N�����d�n�u�u�#�-�B؁�����9��R��]���
�d�3�
�f�d�����ƭ�l��D�����f������1���s���G��V�� ��c�
�d�i�w�)�(�������P������� �&�2�0��?��������U��[�����d�|�n�u�w�)���&����P��N�U���
�:�<�
�2�)�ǫ�
����WN��G]�*���!�6�&�
�"�j�O���P����]��Y������d�3�
�o��E���s���G��1��*��g�%�u�h�u�� ���Yۓ��Z��SF��*���
� �d�`��n�W�������V��G1�����9�d�
�m�~�8����I��ƹF��Z��E���
�e�
�g�k�}�F������@��R
�����d�3�
�m��o�W���������T�����d�
�c�|�2�.�W��B�����hX�����g�
�d�i�w�)�(�������P������� �&�2�0��2�F�������U��Z��D���a�|�_�u�w�0�(�������9��R�����9�2�6�#�4�2�_�������T��D�����4�
�
�
�"�h�C���Pߒ��Z��P�� ���2�0�}�e�w�}����H����T��G_��D��1�"�!�u�~�t�^�ԜY�Ƹ�C9��h��D��
�f�i�u��<�E�������U��F�U���;�:�g�|�]�}�W���&�ғ�F9��1��U��w�w�"�0�w�.����Q����lW��B1�M���|�i�&�2�2�u��������EW��X��U���0�w�w�_�w�}����L����^��G_��Hʦ�1�9�2�6�!�>����������^	��¥�&�
�
�4�#�;�(��&���R�d��U���u�!�%�c��<����&����CW�
N�����2�6�#�6�8�u����ە��]��C��@؊� �c�e�%�~�n�^��s���G��X�� ��e�
�d�i�w�����K����W��h�D���d�1�"�!�w�t�}���Y����Q��B1�G���u�h�w�w� �8�Wǌ�����e9��Q��Mފ�g�h�4�
�8�.�(���M���V
��L�N���u�!�%�c��2�(���@�ޓ�F�F����
� �m�m�'�}����	����@��A_��\�ߊu�u�8�
�o�;�(��&���F�N�����%�&�
�
�"�j�O���Y�ƭ�l��D�����f�|�0�&�w�m�L���YӒ��lP��Q��B���%�u�h�}�6�:�F�������@9��^_��@���
�b�e�%�w�2�W�������l
��h_����u�8�
�
�"�n�O���Y���D��_��]���
�
� �f�e�-�W���	����@��AX��E���9�0�w�w�]�}�W���&�֓�F9��\��G��u�!�%�f��8�(��NӉ��F��E�����'�2�f�`�~�W�W�������l ��V�*��i�u�<�;�0�l����J����K	��V�����
�#�
�|�]�}�W���&�ԓ�F9��]��F��u�
�4�g�d�;�(��N����U��X����|�_�u�u�:��D���&����l��S��D���=�;�}�<�9�9��������l��h]�G���u�<�;�1�6�����&����lV������w�_�u�u�:��C���&����l��S�����:�<�
�0�#�/�����ι�@��R
�����&�2�
�
�"�o�G܁�K����O��N�����b�
� �g�e��E��Yۈ��@��U��G���
�g�l�%�w�2�W�������l
��h_����u�8�
�c�1��E���	���N��P �����2�f�b�u�8�}��������EW��UךU���8�
�b�3��n�E���Y���D��_��]���;�1�%��;��F���&����l��P�����1�4�
�:�$�����I����_��^�����u�8�
�m�1��C���	���N��X������!��0�#�/�8�������@9��h\�M���u�u�:�9�/��8���>����V��E1�� ���d�3�
�f�a�-�^�������K!��x��2���!�'��
�&�<�(�������9��UךU���8�
�l�3��i�C���Y���D��_��]���
�m�3�
�c�i����Y����\��h��*���0�&�u�e�l�}�WϪ�	�ѓ�F9��V��D��u�!�
�:�>�����۔��Z��B �����}�=�4�!�4�.�(���H����CW�Z��N���u�!�%�m��(�E��&���F�N�����!�%�b�
�"�o�Gہ�M����C9��Y�����c�u�9�0�u��}���Y����W��B1�E���u�h�!�%�e����M����W��X����n�u�u�!�'�e�(���K����CT�
N��Wʢ�0�u�!�%�`����Iǹ��[��G1�����9�f�b�u�;�8�U���s���F�C��Mي� �g�b�
�f�a�W���&����P9��T��]���<�0�&�2�2�u�(���K�ޓ�F9��_��F���c�|�_�u�w�}�WϪ�	����U��Y�����h�&�1�9�0�>�����ξ�@�������%��9�
��(�E��&���P�dךU���u�u�8�
�b�;�(��M����[��C
�����
�0�!�'�%�.����������V��@��
� �g�l��n�[��P��ƹF�N�����c�3�
�c�o�-�W��
����\��h�����'�&�/�}�>�3�Ǯ�/����^��B1�@ӊ�f�y�c�|�]�}�W���YӒ��l^��Q��B���%�u�h�&�3�1��������AN��D��]���;�1�<�
�2�4���U���lǻN�����
� �d�l��o�K�������T��A�����=�3�
�<�?�u����ۋ��l0��B1�Fӊ�f�y�:�<�#�:�ǫ�
����WN�N�����b�3�
�e�o�-�_��Hӂ��]��G��\��u�u�!�%�n����@����Z�D�����6�#�6�:��8��������]��F�����;�b�3�
�o�e����J���9F���*���3�
�l�e�'�}�J�������]��h]�� ��e�
�f�-�%�<�(���
����9��d��Uʡ�%�l�
� �e�i�(��E����^��_�����d�g�-�'�6�����&����O��N�����l�
� �g�o��E��Yە��]��h_�����e�d�-�'�6�����&����O��N�����l�
� �f�`��F��Y����_	��T1�����}�0�<�0�"�.����Q����@��Y1�����e�b�%�|�d�t�L���YӒ��l_��Q��E���%�u�h�}�2�.�����ғ�F9��_��Fʭ�'�4�
�:�$��ށ�P���F��G1�*���f�g�
�g�k�}����H�ޓ�V��Z����4�
�:�&��+�(���s���G��Y�� ��c�
�g�i�w�.�����ԓ�V��_����4�
�:�&��+�(���s���G��V�� ��a�
�a�i�w�����&����lW��h��F��
�g�f�u�8�3���B�����hW�����g�l�%�u�j��Uϩ�����q9��h-�����'�6� �0�f�e����M����F��h�����#�
�|�0�$�}�G��Y����^��h��D��
�g�i�u�#�����&����\��Y������
�0�
�`�m�W�������V��G1�����9�d�
��~�f�W�������F9��\��F��u�4�
�:�$��ށ�Y�Ƹ�C9��h��*��b�n�u�u�#�-����&����l��S�����:�<�
�0�#�/��������R��X ��*���g�d�|�x�"�.����Q�ԓ�V�� V�\�ߊu�u��6��<��������A��V�� ��c�
�f�i�w�}�W���Yӕ��l��Y�� ��`�
�f�"�2�}��������F9��W��G��u�u�d�|�2�.�W���Y�����h��@܊� �g�a�
�d�W�W�������lT��1��U��w�w�"�0�w�(�����Ϊ�C9��d�����&�9�!�
�6�(�(���H����T��h�U���;�<�;�1�1�-�6���6����Q��B��#���0�l�
�
�"�o�Oہ�J����_��^�����u�;�0�3�8��(���H����CT�
N�����4�&�2�
��(�F��&����]��E����
�d�3�
�o�d����s���F��E�����3�
�f�a�'�}�J�������l��X�����
�f�m�%�w�2�W�������A��W�\�ߊu�u�;�0�1�2�(݁�����lT��1��U��}�8�d�
�"�o�Eځ�KӉ��C9��h�� ��m�
�g�n�w�}��������lU��B1�Dڊ�g�i�u�&�0�?��������Q��V �����a�3�
�e�c�-�^�ԜY�ƹ�W��[��F���!�3�
�e�`�-�W��Q����9��h]�D���u�'�%�f��l����@�Փ�O��N�� ���'�9�"�a�1��F���	���N��P �����'�2�a�d�w�3�W���HŹ��lU��1��\�ߊu�u�;�0�1�2�(ہ�����lU��1��U��}�8�d�
�"�n�G߁�KӉ��C9��h�����d�g�%�|�]�}�W�������D9��h_�F���u�h�}�<�9�<����&����
T��G]�����'�0�2�l�����OĹ��]��Y
�����n�