-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ���d���}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e�'�3�4�'�<�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y����C9��T��;ʆ�����]�}�W���&����R
��V1��*���u�u�����0���s���C9��E�����o��u����>���<����N��
�����e�n�u�u�'�l��������C9��SN�<����
���l�}�WϮ�K����Z	��N��U���
���
��	�%���Hӂ��]��G�U���%�g��'�8���������}F��s1��2���_�u�u�
����������\��b:��!�����
����_������\F��d��Uʥ�a��!�8�9��(߁�	����\��b:��!�����n�u�w�-�C�������T9��N�:���������4���Y����W	��C��\�ߊu�u�
�
��4�����ד�C9��SN�:��������W�W���&ƹ��U9��C��U���������4���Y����W	��C��\�ߊu�u�
�
�2���������WF��~ ��!�����n�u�w�-�A�������T9��N�:���������4���Y����W	��C��\�ߊu�u�
�
��4�����֓�C9��SN�:��������W�W���&Ź��G��Y	��*���u� �u����>���<����N��
�����e�n�u�u�'�k�5�������V9��V�����u� �u����>��Y����l^��h:�����0�e�o����3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���&����^��h��*���#�1�o����3���>����F�G1��6���8�;�
�
�w�}�"���-����t/��a+��:���f�u�:�;�8�m�L���YӖ��l%��^�����d�4�
�9�w�}�"���-����t/��=N��U���`��6�:�w�}�"���-����t/��a+��:���b�1�"�!�w�t�}���Y����l5��C�����9�u�u� �w�	�(���0���9��dװ���<�0�!�'�w�8����Ӌ��q$��t(��Eʼ�u�u�u�4�#�4����:����t#��e/��:�����o����L���YӇ��A��C��:���������9����Ʈ�[��N�����0�!�'�u�$�}�W���O����%��h^�����%�g�d�
�{��$���)����j6��T��=��������	�FÖ�*����f2��~6��H����
�� ���#Ҧ�N����P
��Z��Y���
�� �
���J��I����J��d1��%�����h�!�2�.�?���*����)��
\�M��e�y��
���6��N߮��l5��h:��H���0������:��1����j(��d>��EƝ�����j�j�OÖ�*����l*��
_�Fި�n�u�u�6�9�)����	����@��X	��*���u��
���}�J���^���F��Y�����%�6�;�!�;�:���Cӵ��l*��~-��H��r�_�u�u�8�.��������l��h��*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-�$�������^9��N��1��������}�E�������V�S��E��e�e�e�e�g�m�G��I���9F������!�4�
��$�n����K����g"��x)��*�����}�g�3�*����P���V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����
�!�
�&��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�n�w�}��������R��c1��@���8�a�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��_�E���_�u�u�:�$�<�Ͽ�&����GP��D��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'��(���&����F��d:��9�������w�o�W������F��L�E��e�e�e�e�g�l�G��I��ƹF��X �����4�
��&�o�;���Cӵ��l*��~-��0����}�g�1� �)�W���C���V��^�E��e�d�e�e�g��}���Y����G����&���!�
�&�
�w�}�#���6����e#��x<��G���:�;�:�e�w�`�U��I����V��^�E��e�e�n�u�w�>�����ƭ�l5��D�*���
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��u�u�6�;�#�3�W���*����W��D��E��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6��#���H����^9��T��!�����
����_������\F��T��W��e�e�e�e�f�m�G��I����l�N�����;�u�%���)�D�������	F��s1��2������u�e�}�������	[�^�E��e�d�e�e�g�m�G��B�����D��ʴ�
��&�d��.�(��Cӵ��l*��~-��0����}�g�1� �)�W���C���V��^�D��e�e�e�e�g��}���Y����G����&���!�`�3�8�f�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�n�w�}��������R��c1��D܊�&�
�`�o���;���:����g)��\����!�u�|�o�w�m�G��I����V��^�E��w�_�u�u�8�.��������l�� 1����u�u��
���(���-���T��X����u�h�w�e�g�m�G��I����V��^�N���u�6�;�!�9�}����&����l ��h_�Oʆ�������8���K�ƨ�D��^��O���e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��	���&����^�=��*����
����u�EϺ�����O�
N��E��e�e�e�e�g�m�G��I����F�T�����u�%��
�#�m����H����`2��{!��6�����u�g�w�2����I����D��_�E��e�e�e�e�g�m�G��Y����\��V ������&�g�
�$��G��*����|!��h8��!���}�g�1�"�#�}�^��Y����V��^�E��e�e�e�e�u�W�W�������]��G1��*���g�3�8�g�w�}�#���6����e#��x<��G���:�;�:�e�w�`�U��I����V��^�E��e�e�n�u�w�>�����ƭ�l5��D�*���
�g�o����0���/����aF�N�����u�|�o�u�f�m�G��I����V��^�E���_�u�u�:�$�<�Ͽ�&����G9��\��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[��D��������4���Y����\��XN�U��w�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��e�d�w�_�w�}��������C9��Y����
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�d�e�w�]�}�W���
������T�����f�
�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�e�d�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�d�g��}���Y����G�������!�9�f�
�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�f�m�U�ԜY�Ư�]��Y�����;�!�9�f��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�l�F���s���P	��C��U���6�;�!�9�d��W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�F��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��H����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��H����l�N�����;�u�%�6�9�)���&���5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��2�����ԓ�F��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-��������9��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��N�&���������W������\F��T��W���_�u�u�:�$�<�Ͽ�&����G9��\��@��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V��^�D��d�n�u�u�4�3����Y����\��h��*���u��
����2���+����W	��C��\��u�e�w�_�w�}��������C9��Y����
�a�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�d�d�e�l�}�WϽ�����GF��h�����#�a�e�o���;���:����g)��X����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�u�W�W�������]��G1�����9�c�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�f�f�W�������R��V�����
�#�g�d�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�c��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��Y����\��V �����:�&�
�#�e�l�W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��H����F�T�����u�%�6�;�#�1�D݁�?�Տ�V�=��*����
����u�FϺ�����O�
N��E��d�d�e�d�g�l�F��H����V��^�����u�:�&�4�#�<�(���
���� T��^�E��o������!���6���F��@ ��U���o�u�d�e�g�m�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D�����d�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�d�w�]�}�W���
������T�����f�
��o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�d�d�g�f�W�������R��V�����
�#�
��m��3���>����v%��eN��U���;�:�e�u�j��F��H���9F������!�4�
�:�$�����I����g"��x)��*�����}�g�3�*����P���V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�f�b�g�$���5����l0��c!��]���:�;�:�e�w�`�U��[���F��Y�����%�6�;�!�;�n�A��*����|!��h8��!���}�u�:�;�8�m�W��[����l�N�����;�u�%�6�9�)����N����g"��x)��*�����}�u�8�3���Y���W��d��Uʶ�;�!�;�u�'�>�����Փ�\��c*��:���
�����}�������	[�^�N���u�6�;�!�9�}��������EU��T��!�����
����_�������V�S��D��n�u�u�6�9�)����	����@��A]��U����
�����#���Q�ƨ�D��^��O���e�e�n�u�w�>�����ƭ�l��D��ي�u�u��
���(���-���F��@ ��U���o�u�e�d�l�}�WϽ�����GF��h�����#�g�f�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�d�d�f��}���Y����G�������!�9�f�
�c�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�f�l�G��Y����\��V �����:�&�
�#�e�n�W���-����t/��a+��:���f�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�l�F��[���F��Y�����%�6�;�!�;�k�(���Y����)��t1��6���u�c�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�l�(��Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���W��^�E��w�_�u�u�8�.��������]��[�*��u�u��
���(���-���V��X����u�h�w�e�g�l�G��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�Fށ�Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��n�u�u�6�9�)����	����@��A_��3���o������!���6���F��@ ��U���o�u�d�d�f�l�F��[���F��Y�����%�6�;�!�;�l�(��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��_�D��n�u�u�6�9�)����	����@��AX��U����
�����#���Q�ƨ�D��^��O���e�e�e�w�]�}�W���
������T�����c�f�u�u���8���&����|4�N�����u�|�o�u�f�m�F���s���P	��C��U���6�;�!�9�b��W���-����t/��a+��:���`�u�:�;�8�m�W��[����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�n�w�}��������R��X ��*���g���o���;���:����g)��_����!�u�|�o�w�l�F��H����D��N�����!�;�u�%�4�3����Lǹ��u ��q(��3���u�u��
���(���-���U��X����u�h�w�d�f�l�F��H����W��_�D��d�d�d�d�f�l�F��H����W��L�U���6�;�!�;�w�-��������9��N��1��������}�F�������V�S��E��e�e�e�e�u�W�W�������]��G1�����9�d�
�c�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����W��d��Uʶ�;�!�;�u�'�>��������F��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-��������lV�=��*����
����u�W������F��L�E��e�n�u�u�4�3����Y����\��h��G������u�w�	�(���0����p2��F�U���;�:�e�u�j��F��H����W��_�D��d�d�d�d�f��}���Y����G�������!�9�f�
��g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�f�l�F��Y����\��V �����:�&�
�#�e�o�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�W�ߊu�u�:�&�6�)��������_��h\�Oʆ�������8���H�ƨ�D��^��O���e�e�e�d�g�m�U�ԜY�Ư�]��Y�����;�!�9�g�d�g�$���5����l0��c!��]���:�;�:�e�w�`�U��B�����D��ʴ�
�:�&�
�!��W���-����t/��a+��:���d�1�"�!�w�t�M���I����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>�����ӓ�\��c*��:���
�����}�������	[�^�E��u�u�6�;�#�3�W�������l
��h]��U���
���
��	�%���Y����G	�N�U��e�d�n�_�w�}����Ӈ��p5��D��U���
���
��	�%���Kӂ��]��G��H���e�e�e�e�g�m�G��I����D��N�����<� �0�3�:�8��������@��Y	�U���4�!�<� �2�;��������TF����6���&�u�u�<�9�1��������l�N�����u�%�&�2�4�8�(���
�ד�@��T��!�����n�u�w�.����Y����Z��S
��L������]�}�W�������lV��R�����
�;�&�2�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������lV��R�����
�'�2�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�f�W���
����_F��1�����%�4�4�
�;���������g"��x)��N���u�&�2�4�w��(���&����R9��h��*���2�o�����4��Y���9F������%�d�'�3�:�%��������`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�d�'�3�8�/�-����Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����F�D�����
�
�0�
�6���������@��N��1�����_�u�w�4����	�ד�V ��V�����1�%�0�u�w�	�(���0����A��d��Uʦ�2�4�u�
��8��������TF��d:��9�������w�n�W������]ǻN�����9�%�g��%�2�(�������g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����9�%�g��%�2�(�������]9��PN�&������_�w�}����Ӗ��l6��^�����9�
�'�2�m��3���>���F�UךU���<�;�9�%�b�/��������l��T��!�����
����_������\F��d��Uʦ�2�4�u�
��8�(�������TF��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���&�2�4�u����������C9��S1��*���u�u��
���L���Yӕ��]��G1�����7�!�
�%�!�9����Y�Ɵ�w9��p'��O���e�n�u�u�$�:��������lR��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�%�:�C��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����2�6�0�
��.�O������5��h"��<��u�u�&�2�6�}��������lW��T��:����n�u�u�$�:����	����l��F1��*���a�3�8�d�w�}�#���6����9F������4�
�<�
�3��F���Y����v'��=N��U���;�9�4�
�>�����J����q)��r/�����u�<�;�9�0�-����H����\��c*��:���
�����l��������l�N�����u��6�
�6�8�$�������lU��1����b�u�u����>���<����N��
�����e�n�u�u�$�:����	����l��F1��*���
�&�
�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�1��i�W���6����}]ǻN�����9�2�%�3��l�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��&����,� �
�f�����N���5��h"��<������}�f�9� ���Y����F�D������6�
�4�2���������9��hZ�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������V9��E�� ���b�
�0�
�`�i�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��G1�����0�
��&�n�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}����&����T��N�&���������W������\F��d��Uʦ�2�4�u�8������A���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�d�
� �b�j����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���'�2�g�e�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������`9��d�����&�9�!�
�6�(�(�������9��T��!�����
����_������\F��d��Uʦ�2�4�u����8���8����F��a����
�0�
�m�e�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������[1��0���!��0�!�%��(�������U��_��G��������4���Y����\��XN�N���u�&�2�4�w�2����<����l!��V��*���� �9�&�%�:�E��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�f�3�
�n��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����
�0�
�m�g�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����R��^	������
�!�e�1�0�N��*����|!��d��Uʦ�2�4�u�%�$�:����H���$��{+��N���u�&�2�4�w���������G��C��*���a�3�
�l��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��d1��*���0��'�6�"�8�Dށ�&����^��T��!�����
����_������\F��d��Uʦ�2�4�u��4�����*����G��h[��F���
�g�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������`9��h-�����'�6� �0�b��(���&����\��c*��:���
�����l��������l�N�����u��6�
�6�8�$�������lR��1��*��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������l%��R1����� �0�a�
��8�(��N����g"��x)��*�����}�d�3�*����P���F��P ��U���6�
�4�0��/�������� 9��hV�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������V9��E�� ���f�
�
�0��e�E��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������4�0��'�4�(���O����
T��G]��U���
���
��	�%���Y����G	�UךU���<�;�9� ��.�4���&����P��R1�C���2�g�`�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӈ��@��T��*���&�d�
�&��l�Mύ�=����z%��N�����4�u�%�&�0�?���@����|)��v �U���&�2�4�u�%����M����	F��s1��2������u�d�}�������9F������3�
�:�0�#�/�(��&����^��T��!�����
����_������\F��d��Uʦ�2�4�u�%�$�:����&����GW��Q��D���u��
���f�W���
����_F��h��*���
�e�u�u���6��Y����Z��[N�����
�l�
�g�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������`9��s*�� ���1�
�e�
�2��O��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V����� �f�l�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����U5��v*��:����1�d�l�%�:�E��Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�������,� ��(���� ����l ��^�����u��
����2���+������Y��E��u�u�&�2�6�}�$���,����F��B�����d�`�'�2�e�e�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��^�����2�g�l�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӈ��@��T��*���&�d�
�&��i�Mύ�=����z%��N�����4�u�%�&�0�?���L����|)��v �U���&�2�4�u�:��D���&����CW�=��*����
����u�FϺ�����O��N�����4�u�8�
�d�/���I����`2��{!��6�����u�`�w�2����I��ƹF��^	��ʡ�%�d�
� �n�j����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���'�2�g�e�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������9��hW�*��o������!���6���F��@ ��U���_�u�u�<�9�1�1݁�����U�=��*����
����u�FϺ�����O��N�����4�u�8�
�b�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�d�
�0��d�C��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��^��D���
�l�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƥ�^��E��G��u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����Aǹ��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Oہ����� P�=��*����
����u�W������]ǻN�����9�<�;�2�f�;�(��@����	F��s1��2������u�g�9� ���Y����F�D�����&�0�
�
�2��N��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����c�3�
�e�d�-�W���-����t/��a+��:���`�u�:�;�8�m�L���Yӕ��]��Z��#���'�2�g�`�w�}�#���6����e#��x<��@���:�;�:�e�l�}�Wϭ�����G��_�� ��l�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����W��R	��L��o������!���6�����Y��E��u�u�&�2�6�}�E�������
Q��N�&���������W��Y����G	�UךU���<�;�9�������@���5��h"��<������}�f�9� ���Y����F�D�����8�
�c�3��l�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����c�'�2�g�`�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h_�*���d�e�
�d�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������^��_�����l�d�o����0���/����aF�N�����u�|�_�u�w�4��������R��B1�Gي�f�o�����4���:����V��X����n�u�u�&�0�<�W���&����A��W�U����
�����#���Q�ƨ�D��^����u�<�;�9�%�l����K�ӓ�F��d:��9�������w�m��������l�N�����u�
�
�0��d�E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��G1��؊�
� �d�l��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��h8��G���'�2�g�l�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����R��^	������
�!�c�1�0�F���Y����)��tUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�)���&����S��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�n�(���&����\��c*��:���
�����}�������9F������1�9�!�1�-�/����&����l��N��1��������}�GϺ�����O��N�����4�u�0�0�2�����&���� V��T��!�����
����_�������V�=N��U���;�9��;�2���������l��1��*��d�%�u�u���8���&����|4�N�����u�|�_�u�w�4����+����9��[1�����
�
�d�'�0�n�F���Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���g�
� �d�a��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����c�'�2�f�f�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������1��*��f�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������A��^�U����
�����#���Q�ƨ�D��^����u�<�;�9�'��݁�I����_��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�'��݁�I����lU��N�&���������W��Y����G	�UךU���<�;�9� �3�/����H����T��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�9�8����&¹��T9��Z��U���
���
��	�%���Y����G	�UךU���<�;�9�%�n���������9��h\�D���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1���&����A��h�����f�a�u�u���8���&����|4�N�����u�|�_�u�w�4��������l%��R1����� �0�d�l�1��A���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʠ�
�!��&��)��������
9��P1�A���u��
����2���+������Y��E��u�u�&�2�6�}��������B9��h��B���8�d�u�u���8���B�����Y�����<�
�1�
�o�}�W���5����9F������ �
�!��$���������Q��Q��C���%�u�u����>���<����N��
�����e�n�u�u�$�:����5����p��h=�� ���'�
�b�
�2��G��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��7���
�4�0��%�>����H�Г�R��Q��C���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϫ�&����R��d�����0�d�c�6�$�����I���5��h"��<������}�w�2����I��ƹF��^	��ʴ�
�<�
�&�&��(���@����lW��N��1�����_�u�w�4��������T9��S1�D������]�}�W�������9��h(��*���%�d�a�3��k�N���Y�Ɵ�w9��p'��#����u�d�1� �)�W���s���@��V��9���
�:�
�:�'�l�C�������F��d:��9�������w�l��������l�N�����u�%�&�2�4�8�(���
����U��W��U���
���n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��G1�*���g�l�
�d�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������^��1����c�u�u����>���<����N��
�����e�n�u�u�$�:��������]��B1�Mي�g�o�����4���:����V��X����n�u�u�&�0�<�W���I����l��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�;��(��&����_	��h��*��e�o�����4���:����U��S�����|�_�u�u�>�3�Ͽ�&����P��h=����
�&�
�d�m��3���>����F�D�����%�&�2�7�3�n�B��;����r(��N�����4�u�!�e�c�h��������`2��{!��6�����u�f�w�2����I��ƹF��^	��ʶ�
�����8���O����l��h]�@��������4���Y����W	��C��\�ߊu�u�<�;�;�?����H����R��R��U����
�����#���Q�ƨ�D��^����u�<�;�9�5�;�G��Mʹ��F��d:��9����_�u�u�>�3�ϼ��֓�R��F^��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�"��(��@����A��N�&���������W������\F��d��Uʦ�2�4�u� ���E������5��h"��<��u�u�&�2�6�}����&����l��T��!�����n�u�w�.����Y����9��W��D��������4���Y����W	��C��\�ߊu�u�<�;�;�?����H����BW�=��*����
����u�FϺ�����O��N�����4�u�!�e�c�h��������@��N��1��������}�FϺ�����O��N�����4�u�!�e�c�h�������5��h"��<��u�u�&�2�6�}����M�ӓ�lV��S
����o������!���6�����Y��E��u�u�&�2�6�}����M�ӓ�lV��R_��U���
���n�w�}�����Ơ�lV��[��*ڊ�0�u�u����>��Y����Z��[N��*ڊ�a�
�
�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W�������
��1�@���e�$�u�u���8���&����|4�^�����:�e�n�u�w�.����Y����lR��h��*���'�&�e�o���;���:����g)��_�����:�e�n�u�w�.����Y����lR��h��*���u�u��
���L���Yӕ��]��[��*��
�
�
�1�%�.�F��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��[��*��
�
�
�0�w�}�#���6����9F������9�
�
�a���(���Y�Ɵ�w9��p'�����u�<�;�9�;��(��&����WW�=��*����
����u�FϺ�����O��N�����4�u�!�e�c�h��������`2��{!��6�����u�f�w�2����I��ƹF��^	��ʼ�
�<��'��2�(������� F��d:��9�������w�l��������l�N�����u�%�&�2�4�8�(���
����U��^��U���
���n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��h��*���$��
�!�o�;���Y�Ɵ�w9��p'�����u�<�;�9�6���������F��u!��0���_�u�u�<�9�1��������V��c1��Gي�&�
�g�o���;���:���F��P ��U���&�2�7�1�c�j�MϜ�6����l�N�����u��6�
�6�8�$�������lW��h��G��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������f*��Y!��*��� �g�d�
�c�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h��F���%�u�u����>���<����N��
�����e�n�u�u�$�:��������lU��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�6�����
����g9��_�����e�o�����4�ԜY�ƿ�T�������7�1�a�l�m��8���7���F��P ��U���
� �f�l�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���M�Փ�F��d:��9�������w�n�W������]ǻN�����9�3�
���$��������_��[�� ��m�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����~3��N!��*���!�%�,�d�b�;�(��&���5��h"��<������}�f�9� ���Y����F�D�����'�
� �a�e�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����d�
�d�o���;���:����g)��]����!�u�|�_�w�}����Ӂ��l ��_�����u��
����2���+������Y��E��u�u�&�2�6�}��������l��N��1��������}�D�������V�=N��U���;�9�2�%�1��Eہ�I����g"��x)��*�����}�f�3�*����P���F��P ��U���&�<�;�3��o�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*���<�;�d�3��n�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V����� �a�f�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����T��Q��Fي�d�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����U��G^��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%����A����	F��s1��2������u�d�}�������9F������!�%�a�
�"�i�D���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����!��&�
�#�(����&�ѓ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(������� 9��T��!�����
����_������\F��d��Uʦ�2�4�u����8���8����F��a����
�
� �`�c�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����a�
�e�o���;���:����g)��^�����:�e�n�u�w�.����Y����U��]��G��������4���Y����\��XN�N���u�&�2�4�w�/�(���M�ԓ�F��d:��9�������w�m��������l�N�����u�'�
� �c�e����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������4�0��'�4�(���&����]��B1�F���u�u��
���(���-��� W��X����n�u�u�&�0�<�W�������@��C�����
�g�;�2�1��Aف�K����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
� �a�a�-�W���-����t/��a+��:���b�1�"�!�w�t�}���Y����R
��Z��*���a�c�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƣ�G��h��A���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϰ�����U��^��G��������4���Y����\��XN�N���u�&�2�4�w�/�(���M�ѓ�F��d:��9�������w�m��������l�N�����u��6�
�6�8�$�������lS��C����� �`�b�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����G��\�� ���d�%�u�u���8���&����|4� N�����u�|�_�u�w�4��������9��h[�*��o������!���6���F��@ ��U���_�u�u�<�9�1�����ԓ�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�9�)��������9��T��!�����
����_�������V�=N��U���;�9�3�
��%��������G��V��*���;�3�
�`��o�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�� ��g�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������l%��R1����� �0�g�
�8�4����&����CW�=��*����
����u�FϺ�����O��N�����4�u��������
����V9��[��G���
� �`�d�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�*���`�b�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lT��Q��M݊�d�o�����4���:����T��S�����|�_�u�u�>�3�ϰ�����l ��_�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�3����M����V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�n�(���L�ӓ�F��d:��9�������w�j��������l�N�����u�8�
�a�1��Gځ�H����g"��x)��*�����}�g�3�*����P���F��P ��U���'�&�
� �a�n����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�� �����
� �c�b�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h]�����g�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����W��B1�L���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����M����lP��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��A���&����CT�=��*����
����u�W������]ǻN�����9�!�%�`��(�A���	����`2��{!��6�����u�d�3�*����P���F��P ��U���
�e�3�
�b��C��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��C���
�l�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƥ�^��B1�F���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������V9��E�� ���f�
� �b�e�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��E�����b�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����G��h��B���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����9��hY�*��o������!���6�����Y��E��u�u�&�2�6�}�$���&����l5��B�����d�c�3�
�e��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������!�3�
�`��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�����m�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����G��h��B���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����9��hY�*��o������!���6�����Y��E��u�u�&�2�6�}�$���&����l5��B�����d�b�3�
�c��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���c�1�8�'�6����@����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�d��8��������Q��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�i����@ù��\��c*��:���
�����}�������9F������&�9�!�%�1��Oځ�K����g"��x)��*�����}�u�8�3���B�����Y�����!��&�
�#�(����&�ד�l �� Y�����u��
����2���+������Y��E��u�u�&�2�6�}�$���&����l5��B�����g�d�3�
�g��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������4�0��'�4�(���&����l^��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�1�����
����A��B��@؊� �b�m�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����@��C��*���m�m�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƿ�_9��GW�� ��`�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G��h��M���%�u�u����>���<����N��
�����e�n�u�u�$�:����*����p��h=�� ���'�
�m�3��h�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��&���
�4�0��%�>����J˹��U��]��F��������4���Y����W	��C��\�ߊu�u�<�;�;�;�(���:����`��T����
�
� �m�f�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��C��@ފ� �m�f�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�����m�
�f�o���;���:����g)��\�����:�e�n�u�w�.����Y����G9��D�����!�'�
�
�"�j�B���Y�Ɵ�w9��p'��#����u�g�1� �)�W���s���@��V�����b�3�
�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�e�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��E���
�l�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƨ�R��P �� ��b�%�u�u���8���&����|4�]�����:�e�n�u�w�.����Y����l0��B1�F���u�u��
���(���-���U��X����n�u�u�&�0�<�W���&����e9��hW�*��o������!���6���F��@ ��U���_�u�u�<�9�1����Lʹ��l_��h�Oʆ�������8���O�ƨ�D��^����u�<�;�9�#�-����&����CW�=��*����
����u�FϺ�����O��N�����4�u�8�
�n�;�(��&���5��h"��<������}�g�9� ���Y����F�D�����8�
�l�3��m�F���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����m�
� �d�f��F��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��Fڊ� �d�e�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����C9��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:����&����T��h��A���%�u�u����>���<����N��
�����e�n�u�u�$�:��������lW��B1�Fۊ�d�o�����4���:����P��S�����|�_�u�u�>�3�ϻ�	����l0��h��D��
�a�o����0���/����aF�N�����u�|�_�u�w�4��������V��B1�Cۊ�d�o�����4���:����S��S�����|�_�u�u�>�3�Ϫ�	����U��X�����u��
����2���+������Y��E��u�u�&�2�6�}�(�������l ��^�*��o������!���6��� F��@ ��U���_�u�u�<�9�1����/�Փ�F9�� Y��G��������4���Y����W	��C��\�ߊu�u�<�;�;�)���A����V��h�Oʆ�������8���O�ƨ�D��^����u�<�;�9�#�-�Cց�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��k����H�Փ�F��d:��9�������w�l�W������]ǻN�����9�!�%�c��<����&����l��N��1��������}�D�������V�=N��U���;�9�!�%�f�h����H�ד�F��d:��9�������w�l�W������]ǻN�����9�!�%�c��(�F��&���5��h"��<������}�f�9� ���Y����F�D�����8�
�d�
�"�l�Bց�H����g"��x)��*�����}�u�8�3���B�����Y�����b�
� �d�b��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��G1��D���
�d�f�%�w�}�#���6����e#��x<��@ʱ�"�!�u�|�]�}�W�������^��Y�� ��c�
�f�o���;���:����g)��[�����:�e�n�u�w�.����Y����W��Q��D���%�u�u����>���<����N��
�����e�n�u�u�$�:��������
9��h_�D���u�u��
���(���-���U��X����n�u�u�&�0�<�W���&����U��V�����u��
����2���+������Y��E��u�u�&�2�6�}�(�������l ��_�*��o������!���6��� F��@ ��U���_�u�u�<�9�1����J����W��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�:��E���&����l��N��1��������}�GϺ�����O��N�����4�u�8�
�b�;�(��H����	F��s1��2������u�b�}�������9F������%��&�9�����H˹��\��c*��:���
�����n��������l�N�����u�4�
�
��(�F��&���5��h"��<������}�d�9� ���Y����F�D�����8�
�f�3��o�B���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����a�3�
�g�g�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��q\��*���d�a�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������R��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������
9��h_�C���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1�1݁�&����l ��\�*��o������!���6���F��@ ��U���_�u�u�<�9�1����Kù��lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������P��N�&���������W��Y����G	�UךU���<�;�9�!�'�k�(���H����CW�=��*����
����u�FϺ�����O��N�����4�u�8�
�`�;�(��I����	F��s1��2������u�g�9� ���Y����F�D�����8�
�d�3��o�E���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����9�
�
�
�f�;�(��O����	F��s1��2������u�d�}�������9F������!�%�g�
�"�l�E݁�K����g"��x)��*�����}�d�3�*����P���F��P ��U���
�`�6�&��(�F��&���5��h"��<������}�f�9� ���Y����F�D�����8�
�a�3��n�@���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����c�3�
�f�f�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��L���
�f�c�%�w�}�#���6����e#��x<��@���:�;�:�e�l�}�Wϭ�����G��Z�� ��a�
�g�o���;���:����g)��[����!�u�|�_�w�}����Ӓ��l_��Q��F���%�u�u����>���<����N��
�����e�n�u�u�$�:����&����_��h��D��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������9��h_�B���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������U��^�����u��
����2���+������Y��E��u�u�&�2�6�}����I����lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�%�;�(��J����	F��s1��2������u�g�9� ���Y����F�D�����
�
�
� �f�d�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*���d�f�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƽ�l��^	��D���
�f�c�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��1��*��g�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����_T��h��D��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������U��B1�D؊�f�o�����4���:����V��X����n�u�u�&�0�<�W���&���� 9��h_�F���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l ��Z�*��o������!���6�����Y��E��u�u�&�2�6�}����@����U��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����R��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)��������P��N�&���������W��Y����G	�UךU���<�;�9�&�;�)��������^��N�&���������W������\F��d��Uʦ�2�4�u�0��0�Fׁ�����9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�A���&����l��N��1��������}�D�������V�=N��U���;�9�&�9�#�-�B�������]9��h_�M���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����A����T��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����^��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)��������_��N�&���������W������\F��d��Uʦ�2�4�u�8��n����J�Փ�F��d:��9�������w�n�W������]ǻN�����9�&�9�!�'�d����M�֓� F��d:��9�������w�n�W������]ǻN�����9�!�%�d��2�(���H����CT�=��*����
����u�W������]ǻN�����9�;�!�&�;�)����&����l��N��1��������}�GϺ�����O��N�����4�u�8�
�a�;�(��I����	F��s1��2������u�g�9� ���Y����F�D�����8�
� �d�f��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��G��*���d�g�
�g�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������\��Q��@���%�u�u����>���<����N��
�����e�n�u�u�$�:��������9��h_�L���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����&����l ��[�*��o������!���6���F��@ ��U���_�u�u�<�9�1����Jʹ��lW��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(�������Q��N�&���������W��Y����G	�UךU���<�;�9�9��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʧ�#�
� �d�a��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��*���d�m�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9�� 1��*���l�%�u�u���8���&����|4�N�����u�|�_�u�w�4�������� 9��h_�F���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����&����V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�%�$���������W��N�&���������W��Y����G	�UךU���<�;�9�!�'�i�(���H����CW�=��*����
����u�DϺ�����O��N�����4�u�4�2�e��F���&����l��N��1��������}�B�������V�=N��U���;�9�'��1��A���	����`2��{!��6�����u�`�w�2����I��ƹF��^	��ʺ�
�:�1�d�>�;�(��@����	F��s1��2������u�g�9� ���Y����F�D�����4�2�g�4�;�2��������9��T��!�����
����_�������V�=N��U���;�9��;�2���������l��B1�A݊�f�o�����4���:����V��X����n�u�u�&�0�<�W����ד�_
��Y��D���
�`�f�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��1��*��b�%�u�u���8���&����|4�N�����u�|�_�u�w�4����+����9��[1�����3�
�c�f�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W�������4��P�����/�'�&�d�1��A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�f�;�!�1��@���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�b�3�
�a�h����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���g�
� �d�g��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����f�3�
�b�b�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E1����
�
� �d�b��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��e��ۊ�9�
�;�&�1��A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�g�
�"�l�Eށ�J����g"��x)��*�����}�u�8�3���B�����Y����
�
� �d�n��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��G1�*��� �d�b�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��@���
�b�b�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������R��h_��*���d�g�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƞ�]��h��*���&�g�<�3��j�N���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����d�4�9�/�%�.�E�������S��N�&���������W������\F��d��Uʦ�2�4�u�0�$�:��������S��N�&���������W������\F��d��Uʦ�2�4�u�8��n����N�ߓ�F��d:��9�������w�m��������l�N�����u�8�
�`�1��@���	����`2��{!��6�����u�d�w�2����I��ƹF��^	��ʓ�
�
� �d�o��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*��
� �d�e��i�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h[�����3�
�b�c�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�*���d�g�
�d�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������^��1��*��c�%�u�u���8���&����|4�]�����:�e�n�u�w�.����Y����^��B1�Eڊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����U��]�����u��
����2���+������Y��E��u�u�&�2�6�}�(���K�֓�l��B1�Fߊ�f�o�����4���:����U��S�����|�_�u�u�>�3�Ϫ�	����U��[�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�-�!���&˹��lW�� 1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(��&����Q��G_��U���
���
��	�%���Y����G	�UךU���<�;�9�'�>�4�(���H����CT�=��*����
����u�W������]ǻN�����9�$�
�
�"�l�A߁�J����g"��x)��*�����}�u�8�3���B�����Y�����&�<�;�f�1��O���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�f�3�
�o�d����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��#���
�
� �d�n��E��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*��
� �d�l��n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�l�l�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��Fފ� �d�g�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��\�����m�c�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��[�� ��f�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����G��1��*��f�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G�� 1��*��a�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��h��D���
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CU��Q��L���%�u�u����>���<����N��
�����e�n�u�u�$�:��������CW��h
�����;�3�
�l�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��T��*���d�d�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��GZ�����l�l�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��_�� ��b�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����R��B1�A؊�g�o�����4���:����U��S�����|�_�u�u�>�3�ϭ����� _��B1�@܊�f�o�����4���:����U��S�����|�_�u�u�>�3�Ϫ�	����]	��Q��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϰ�����l��1��*��`�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������9��h_�B���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����&����V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�%�$��(���K����CT�=��*����
����u�FϺ�����O��N�����4�u�:�g�f�;�(��K����	F��s1��2������u�f�}�������9F������!�%�d�c�1��G���	����`2��{!��6�����u�e�3�*����P���F��P ��U���d�d�6�&��(�E��&���5��h"��<������}�f�9� ���Y����F�D�����8�
�b�3��m�N���Y�Ɵ�w9��p'��#����u�`�u�8�3���B�����Y�����b�
� �g�a��E��*����|!��h8��!���}�f�1�"�#�}�^�ԜY�ƿ�T����D���
�e�m�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V��Q��E���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	ƹ��lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�@ځ�����
9��T��!�����
����_�������V�=N��U���;�9�!�%�f�e����I�ғ� F��d:��9�������w�m��������l�N�����u�8�
�e�1��G���	����`2��{!��6�����u�e�3�*����P���F��P ��U���a�3�
�e�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��X��D���&�
� �g�e��F��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T����*���3�
�d�e�'�}�W���&����p9��t:��U���u�:�;�:�g�f�W���
����_F��Y	��*���
� �g�d��o�Mύ�=����z%��r-��'���f�1�"�!�w�t�}���Y����R
��h8��*���g�d�
�g�m��3���>����v%��eN��Fʱ�"�!�u�|�]�}�W�������A9��Y
�*���3�
�d�a�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W�������4��P�����:�0�
�
�"�o�Eځ�K����g"��x)��*�����}�u�8�3���B�����Y��'���0�
�9�
�9�.�F���&����U��G]��U���
���
��	�%���Y����G	�UךU���<�;�9��9�8�(���&����lU��B1�BҊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&�Փ�F9��_��G��������4���Y����\��XN�N���u�&�2�4�w�<��������V��h\�� ��`�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����VW��[�����
�
� �g�`��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��Mڊ�:�
� �g�o��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��Mߊ� �g�c�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��G���
�d�g�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���g�l�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƣ�l��SW��ۊ� �g�f�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����a��R_�����;�&�g�3��l�B���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�a�
� �e�m�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��Lߊ�d�3�
�d�g�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��hW��ۊ� �g�c�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��@���
�g�e�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������R��h_��D���
�e�b�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������R��1�����0�
�
�d�1��E���	����`2��{!��6�����u�e�3�*����P���F��P ��U���2�d�4�9�-�/����¹��lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9��3�ށ�����V��h��D؊� �g�a�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����]��^	�����
� �g�f��n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�g�c�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������1��*��g�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��h��G��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������l ��\�*��o������!���6�����Y��E��u�u�&�2�6�}��������U��X�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)�؁�����9��T��!�����
����_�������V�=N��U���;�9�1�9�#�9����
�ד�F9��X��F��������4���Y����\��XN�N���u�&�2�4�w�8�(���K˹��lT��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Cׁ�����9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�@���&����l��N��1��������}�GϺ�����O��N�����4�u�8�f�1��D���	����`2��{!��6�����u�e�3�*����P���F��P ��U���0�3�:�
�"�o�F߁�J����g"��x)��*�����}�u�8�3���B�����Y����
�0�:�2�9�4����J�ԓ�F��d:��9�������w�m��������l�N�����u�;�0�3�8���������9��T��!�����
����_�������V�=N��U���;�9�%�l��8��������\��B1�Fӊ�g�o�����4���:����V��X����n�u�u�&�0�<�W�������Z9��Y�����f�f�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӓ��lP��Q��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϼ�����l ��]�*��o������!���6�����Y��E��u�u�&�2�6�}��������U��Y�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	�ד�F9�� [��G��������4���Y����\��XN�N���u�&�2�4�w�����H����Z9��O1��*��d�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G��1��*��f�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����A ��@1�����3�
�f�l�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W��������� 1�����4�
�f�f�9�)����J�ߓ�F��d:��9�������w�m��������l�N�����u�'�0�2���D�������F9��Z��G��������4���Y����\��XN�N���u�&�2�4�w�0�(�������Q��N�&���������W������\F��d��Uʦ�2�4�u�'�2�:�F���&����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�h�(���K����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�l����M�Փ�F��d:��9�������w�m��������l�N�����u�
�4�g�f��(��K����l ��Z�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������l ��Z�*��o������!���6���F��@ ��U���_�u�u�<�9�1����J����lT��h�����
� �g�f��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��Z�����a�b�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƹ�l��x��G���9�6�9��1��D���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʠ�
�:�0�!�%��Eׁ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u��4�����*����G��h_�*ۊ� �g�`�
�c�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������T������'�6� �2�l�A�������^��N�&���������W��Y����G	�UךU���<�;�9� ��)�4���&����P��R1�L���3�
�a�g�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�*���g�m�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��h��G��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CS��Q��@���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����_��S�����
� �g�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���g�l�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G[�����`�g�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��^�����'�4�
� �e�n�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
� �g�l��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��[1�����3�
�`�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��@݊� �g�a�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��@���
�`�m�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���g�d�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƹ�l��t��*��� �!�'�
�o��(���K����CT�=��*����
����u�FϺ�����O��N�����4�u�'�6�9����Où��\��c*��:���
�����}�������9F������;�"�0�
�"�o�B݁�J����g"��x)��*�����}�d�3�*����P���F��P ��U����9�
� �e�k�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����;�d�3�
�b�i����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T�������g�3�
�`�b�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R��ي� �g�m�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������d��*���g�m�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������V��[[�� ��e�
�f�o���;���:����g)��]����!�u�|�_�w�}����ӈ��`��h��G��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������_^��B1�F؊�f�o�����4���:����U��S�����|�_�u�u�>�3�ϰ�����l ��X�*��o������!���6���F��@ ��U���_�u�u�<�9�1�����ғ�F9��V��F��������4���Y����W	��C��\�ߊu�u�<�;�;�3� ���Hù��lT��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�8�$���&����S��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�:��B���&����l��N��1��������}�GϺ�����O��N�����4�u��!�%�l�>�������R��t�����
� �g�e��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��{1�� ��� �
�d�
�"�o�F݁�K����g"��x)��*�����}�d�3�*����P���F��P ��U���-� ��;�"��Fځ�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�'��(�D�������`2��{!��6�ߊu�u�<�;�;�:����&����P�=��*����n�u�u�$�:��������lR��h��Oʆ�����]�}�W�������C9��P1������&�g�3�:�l�Mύ�=����z%��N�����4�u�%�&�0�?���J����q)��r/�����u�<�;�9�6�����
����g9��1����o������}���Y����R
��G1�����1�d�a�u�w��;���B�����Y�����<�
�&�$���ہ�
����	F��s1��2���_�u�u�<�9�1��������W9��_��U�����n�u�w�.����Y����Z��D��&���!�
�&�
�w�}�#���6����9F������4�
�<�
�3��A��CӤ��#��d��Uʦ�2�4�u�%�$�:����&����GP��D��U����
���l�}�Wϭ�����R��^	�����c�c�o����9�ԜY�ƿ�T��	��*���a�m�6�u�w�	�(���0��ƹF��^	��ʲ�%�3�
�g��8�Mύ�=����z%��N�����4�u�'�
�"�i�D�������	F��s1��2������u�c�9� ���Y����F�D�����'�
� �a�o�2����Y�Ɵ�w9��p'��#����u�a�1� �)�W���s���@��V�����c�3�
�a��-����Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*���3�8�o����0���/����aF�N�����u�|�_�u�w�4��������T9��S1�U������n�w�}�����ƭ�l��h��*��o�����W�W���������D�����b�u�u����L���Yӕ��]��V�����1�
�m�o���2���s�����G�����c��d��1�m����&�Ԣ�lU��D1�*ي� �9�1�%��W�W�������PF�N��U����u�u����L���Y���(��h=��2���u����l�}�W���Yӂ��9��s:��Oʜ����_�w�}�W����ד�z"��T��;����n�u�u�w�}����&����{F��~ ��2���|�_�u�u�8�)�_���Y�����T��;ʆ�����]�}�W���Y����GF��~ ��!�����n�u�w�}�WϺ�����z(��c*��:���
�����l��������l�N��Uʱ�;�u�u����;���:����g)��]����!�u�|�_�w�}�W�������}F��s1��2���_�u�u�u�w�2���6����g"��x)��*�����}�d�3�*����P����F�R �����:�0�!�_�]�}�W���	����GF��r,��D���
�
�8�9�d�3�(���
����9��O1��ʜ�_�u�u�0�2�4�W�ԜY���F��T��;����n�u�u�w�}�9���*����\��y:��0��u�u�u�u�3�3�(���-����z(��p+�����u�u�u�<�f�
�3���Cӯ��v!��d��U���u�1� �
��	�W���7����aF�=N��U���!�}�u�u�w�}����Y�ƅ�5��h"��<������}�f�9� ���Y����F�N�����u�u�����0���/����aF�N�����u�|�_�u�w�}�W�������f2��c*��:���
�����l��������O��N�����6�8�:�0�#�W�}���Y����\��CN��0���d��
�
�3�+�Dݰ�&�Ԣ�lU�� N�����u�0�0�<�w�W�W���Y�ƅ�\��y:��0��u�u�u�u���$���<����}2��r<�U���u�u�1�;���#���Y����t#��=N��U���u�<�d����Mϗ�-����l�N��Uʱ� �
���w�}�9���<���9F������u�u�u�u�4�6�Mϗ�Y����)��tUךU���u�u�0�0�w�}�9ύ�=����z%��N��U���1�;�u�u���3���>����v%��eN��Dʱ�"�!�u�|�]�}�W���Y����\��yN��1��������}�D�������V�=N��U���u�0�o��w�	�(���0��ƹF�N�����o������0���/����aF�N�����u�|�|�_�w�}��������V��=dךU���:�%�;�;�w�k�5��:����l��X��C޻�
�g�g��]�}�W�������l�N��Uʜ�u�u����f�W���Y����f+��c/��U������n�w�}�W�������d/��N�<�����_�u�w�}�W�������g.�'��0���u�n�u�u�'�/�W�ԜY���F��\N�<����
���l�}�W���YӔ��V�'��&������_�w�}�W������/��d:��9�������w�k�W������]ǻN��U���0�o��u���8���B���F�
����������4���:����U��S�����|�|�_�u�w�3�W���	����G]Ǒ=N��U���%�;�;�u�a��Fޝ��֓�C��h]����
�u��u�w�:������ƹF�N��1������]�}�W���Y����`2��rN�<�����_�u�w�}�W���I����g.�'��0���n�u�u�u�w�9����0����	F��c+��'���_�u�u�:�#�u�W���Y����Z��N��U���
���
��	�%���Hӂ��]��G�U���u�u�1� �w�}�"���-����t/��a+��:���c�u�:�;�8�m�W��Y����]��X�����n�_�u�u�4�0����Ӌ��q$��t(��E���8�
�g�&�d�3�(ށ�Y��ƹF��R �����_�u�u�u�w��Mϗ�-����l�N��Uʛ�����m��#���+���F�N��ڊ���u�u���2��Y���F��^ ��"����o�����}���Y���W	��h9��!���u����w�f�W���	����l�N��Uʱ�;�u�u����;���:����g)��]����!�u�|�_�w�}�W������/��d:��9�������w�n�W������]ǻN��U���%�:�0�o��}�#���6����e#��x<��Aʱ�"�!�u�|�]�}�W���Y����\��b:��!�����
����_�������V�UךU���;�u�:�%�9�3�L�ԶY����\��Y��U����d��3�g�?����H����z5ǻN�����<�u�_�u�w�}�W�������[F��~ ��2���_�u�u�u�w�9����+����\��y:��0��u�u�u�u��9��������	F��c+��'���_�u�u�:�#�u�W���Y����_�'��&������_�w�}�W�������	F��=��*����n�u�u�w�}��������	F��=��*����
����u�W������]ǻN��U���0�u�u����;���:���F�N��U��� �u��
���(���-��� W��X����n�u�u�u�w�<����
����z(��c*��:���
�����}�������9F�N��U���u�u�����0���s���F�@�Oʜ�u��
���f�W���Y����F��~ ��!�����
����_������\F��d��U���u�$�u�u��}�#���6����e#��x<��F���:�;�:�e�w�f�W�������\��Y��N�ߠu�u�6�8�8�8�ϳ�<����p ��1��*ڊ�a�
�
�u��}�WϹ�����NǻN��U���4�4�<�!�w�}�9���<��ƹF�N�����&��;�0�m��#���+���F�N�����&�<�!�u�w��2���Y��ƹF��X��]���u�u�u�6�<�g�>���-����t/��=N��U���u�0�0�u�w��$���5����l�N��Uʴ�1�0�&�u�w��$���5����l0��c!��]���:�;�:�e�l�}�W���YӅ��\��yN��1�����_�u�w�}�W��Cө��5��h"��<������}�g�9� ���Y����F�N�����0�&�u�u���3���>����v%��eN��U���;�:�e�n�w�}�W������/��d:��9����_�u�u�w�}����Y����g"��x)��N���u�u�u�1�w�}�9ύ�=����z%��r-��'���e�1�"�!�w�t�}���Y���BW�!��U���
���
��	�%���Iӂ��]��G��N���u�0�1�6�:�2����s����V��=N��U���
�
�g�l��g����������u,�6���e�7�3�e�f�i�}���Y����A��Z��]���u�u�u��#�
����D����l�N��Uʔ�1�0�&�4�0�}�I��s���F�v
�����<�!�u�k�e�W�W�������R�=N��U���u�9�u�k�6����Y���F��R��U��4�
�&�y�w�}�W�������@��
P�� ���
�g�l�4�3�8���Y���F��R^��Kʷ�3�e�d�a��8�[���Y�����
P�� ���
�g�l�$�{�}�W���YӇ��A��N��U���
�
�g�l�6�9����U���F���U��7�3�e�d�c����Y���F��R_��Kʷ�3�e�d�a��8�[���Y�����
P�� ���
�g�l�1�{�}�W���Yӗ��X��B��*��l�$�|�_�w�}����&����V9��bN����:�0�!�8���F���&ù��lV��[��*�ߊu�u�0�0�>�}����s���F�s��"���=�h�u�d�]�}�W���Y����V��V ��U��f�_�u�u�w�}����
����G�	N����u�:�!�8�'�u�W���Y����_�	N��*���y�u�u�u�w�/����D�ƭ�l��d��U���u�4�1�0�$�}�Iϲ�&ù��9��1�����&�y�u�u�w�}���D�Ơ�lV��[��*ڊ�0�y�u�u�w�}����Gӊ��9��1��E���y�u�u�u�w�<����
���
��1�@���e�4�1�0�$�q�W���Y����VW�	N��*ڊ�a�
�
�
�2�q�W���Y����VW�	N��*ڊ�a�
�
�
�2�q�W���Y����F���E��`�0�e�1�{�}�W���Yӗ��X��C1��A���0�e�$�|�]�}�Wϲ�&ù��9��1��Oʶ�8�:�0�!�:��5���?����Q��1�A�ߊu�u�0�0�>�}����s���F�s��"���=�h�u�g�]�}�W���Y����V��V ��U��f�_�u�u�w�}����
����G�	N����u�:�!�8�'�u�W���Y����_�	N��*���y�u�u�u�w�/����D�ƭ�l��d��U���u�4�1�0�$�}�Iϲ�&ù��9��1�����&�y�u�u�w�}���D�Ơ�lV��[��*ۊ�0�y�u�u�w�}����Gӊ��9��1��D���y�u�u�u�w�<����
���
��1�@���d�4�1�0�$�q�W���Y����VW�	N��*ڊ�a�
�
�
�2�q�W���Y����VW�	N��*ڊ�a�
�
�
�2�q�W���Y����F���E��`�0�d�1�{�}�W���Yӗ��X��C1��A���0�d�$�|�]�}�Wϸ�I����W9��Y��G���f�
�
� �;�9����Y�Ư�^��R ��ܐ��d��
��<�������]��1�����
�&�_�u�w�8����Y����l�N��Uʜ�u�k�d�_�w�}�W���,����r!��
P��Y���u�u�u�1�9��>���Y���JǻN��U���<�d����`�W��s���F�S��*����u�k�f�~�}�WϮ��ơ�CF�N��U���6�>�h�u�'�>��ԜY���F��D��H���%�'�!�_�w�}�W������F��G1��*��
�e�_�u�w�}�W���H���T��Q��Lߊ�d�_�u�u�w�}���Y����U��[���ߊu�u�u�u�8�)�J�������lU��h�N�ߊu�u�
�
�6�9�Dݰ�&�Ԣ�lU��1�����&�
�d�o�4�0����Ӌ��q$��t(��E���1�
�g�&�d�3�(���J����_9��Gd��Uʲ�;�'�6�8�'�u�W���Y����wF�_�U���u�u�����2��Y��ƹF�N��������h�w�o�}���Y���W��h9��!���k�f�y�u�w�}�WϺ�����w2��
P��G�ߊu�u�:�!�:�-�_���Y�����S����9�y�u�u�w�}�������R��D�U���u�u�1�;�w�c��������
9��d��U���u�1�;�u�i�:����&����CW�N��U���6�u�k�2�'�;�(��&����F�N�����u�k�2�%�1��Nց�K��ƓF�Q1�����
�g�&�f�9��E�������@��N����:�0�!�8���F���&ù��F
�� ��Fػ�
�g�d�8�/�9����YӁ��V����U�ߊu�u�u�u��`�W��Y���F��b#��!���u�k�d�_�w�}�W����֓�z"��S�F���u�u�u�u�3�3�(���-���U��=N��U���u�:�!����J���K���F��E�����_�u�u�u�w�4�G��Y����U��]��E�ߊu�u�u�u�>�l�J�������lR��h����u�u�u�:�#�`�W���&����U��G����u�
�
�8�;�n����K����9��Z����� �u�u�:�'�3����O����%��h^�����f�;�
�g�$�n�(ށ�����Cl�N�����6�8�%�}�w�}�W���0���W�N��U��������`�W��Y���F��^ ��"����h�u�g�]�}�W���Y����l1��c&��K��y�u�u�u�w�9����0����X�GךU���:�!�8�%��}�W���Yӂ��F��������!��;�4����Kƹ��lR��h����u�u�u�<�f�`�W�������J)��h#�����,�d�`�3��m�(��s���F�S��U��3�
���.�(�(�������lW��h��A���%�|�_�u�w�;�G�������]�� ��F؊�
�a�o�6�:�2����ţ��W��Q1�����
�g�&�f�9��E��Y����V��^�����_�u�u�u�w��J���U���F� ��*����u�k�b�]�}�W���Y����l1��c&��K��y�u�u�u�w�9�ށ�0����X�BךU���u�u�:�!� ��?��Y���F�G��U���u�_�u�u�w�}����GӇ��P
��=N��U���u�0�0�u�i�<�(���U���F�
��E��u�'�
� �c�o���Y���F��^ �H���'�
� �a�e�-�[���Y�����
P����� �a�g�6�{�}�W���Yӂ��GF�	��*���a�g�%�|�]�}�Wϸ�I����E9��Y��G���f�
�
�`�m�>��������#��_�����3�<�
�g�$�n����K��ƹF��R �����4�u�_�u�w�}�W���D����9F�N��U���
���u�i�j�}���Y���W��h9��!���k�f�y�u�w�}�WϺ�¹��w2��
P��G�ߊu�u�u�u�8�)� ���1��� T�N�����u�4�u�_�w�}�W��������T�����u�u�u�0�2�}�IϿ�&����9F�N��U���e�h�u�'��(�C���	��ƹF�N����h�u�'�
�"�i�O���U���F���H���'�
� �a�o�>�[���Y�����CN��U���
� �a�m�'�t�}���YӀ��l��X��C޻�
�g�g� �w�}��������^P��u_��3���
�<�:�%�a�3�(���K�����R��U���u�_�u�u�w�}�3��Y��ƹF�N�� �����u�k�e�W�W���Y�ƨ�]V��~*��U��c�y�u�u�w�}����&����{F�]����u�:�!�8�'�u�W���Y����_�	N��*���y�u�u�u�w�/����D�ƭ�l��d��U���u�1�;�u�i�:����&����CV�N��U���6�u�k�2�'�;�(��&����F�N�����u�k�2�%�1��Eہ�H��ƓF�Q1�����!�f�;�
�c�l�"���Y����\��CN��0���d��
�
�'�%�(���
����l�N�����6�8�%�}�w�}�W���0���W�N��U��������`�W��Y���F��^ ��"����h�u�g�]�}�W���Y����l1��c&��K��|�u�u�%�%�}����s���F�S��U��1�4�&�2��(�C���	��ƹF�N�����h�u�
�&�>�3����KĹ��]ǑN�����3�0�!�f�9��C���,����P	��X ��ʸ���d�������&�Ԣ�lP��d��Uʲ�;�'�6�8�'�u�W���Y����wF�_�U���u�u�����2��Y��ƹF�N��������h�w�o�}���Y���W	��h9��!���k�c�|�u�w�-�������F�N�����u�k�1�4�$�:�(ށ�����l��=N��U���u�:�!�h�w������ד�F9��1��\�ߠu�u�3�e�1�0�(���
����@9��1��U���:�%�;�;�w�k�5��:����l ��G1����g�&�d�d�w�}��������R�=N��U���u��h�u�{�}�W���YӨ��l5��p+��K��_�u�u�u�w�4�G���=���F��d��U���u�1�;�
��	�W���J��ƹF�N��������h�w�t�W���	����^��d��U���u�1�;�u�i�:����&����CV�N��U���1�;�u�k�0�-����J����l�N��Uʺ�6�1�u�k�0�-����J����P	��d��U���u�1� �u�i�:����&����CT�=d��Uʳ�e�3�8�
�e�.�Dݰ�&¹��fW��N�����0�!�8���l�1���&����lU��D1����
�_�u�u�2�8�������F�N��<���k�d�_�u�w�}�W���&����vF�_�U���u�u�1�;���#���G����9F�N��U���d����j�}�E�ԜY���F��B��<���u�k�d�_�w�}�������9F�N��U���e�h�u�'��(�C���	��ƹF�N����h�u�'�
�"�i�O���U���F������h�u�'�
�"�i�O�������9F�N��U���!�h�u�'��(�C���	����9F���*���%�f�;�
�e�.�F���,�����G�����c��d��1�m����&�Ԣ�lU��D1��D���u�2�;�'�4�0����Y���F��sN��U���u�u�u�u���$���<���JǻN��U���<�e����`�W��s���F�S��*����u�k�f�{�}�W���Yӂ��G9��s:��H���|�u�u�%�%�}����s���F�S��U��!�%�a�
�"�i�D���U���F�
��D��u�8�
�c�1��C܁�H���F�N�����u�k�!�%�c����J����\��=N��U���u�:�!�h�w�0�(������� 9��Uװ�ߠu�u�x�u�?�}�����ƿ�R����6���&�|�:�u�?�}����Y����Z��C�U���4�
��3�:�<����&����\��E�����%�6�>�_�w�}����s���F�^�����9�r�#�;�w�3�W������F�G�����u�u�u�u�w�}��������GF�_��U���;�u�u�u�w�}�W���YӇ��p5��D��Hʴ�
��&�d�1�0�G�ԜY���F�N���ߊu�u�u�u�w�}�W�������C9��Y�����6�d�h�4��8�^Ϫ���ƹF�N��U���u�u�u�u�'��(���Y����C9��h��N���u�u�u�u�w�}�Wϻ�ӏ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���T�Ƽ�9��Q1�����4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�e�'�1�<��������W9��R	�����;�%�:�u�w�/����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�p�z�W������F�N��U���}�%�'�!�j�z�P�����ƹF�N��U���u�u�
�
�2�����&����_��E��I���%�6�;�!�;�:���s���F�N�����_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���K����^9��G�����_�u�u�u�w�}�W���Y���F�G1�����4�%�4�4��1�(������R��X ��*���<�
�n�u�w�}�W���Y���F������4�
�<�
�3��@������F�N��U���u�u�u�u�w�}��������_��h�����%�0�u�h�'�m��������l��A�����u�u�u�u�w�}�W���Y����Z ��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����R
��V1�����&�<�;�%�8�8����T�����h��*���=�
�'�2�6�.���������T��]���6�>�_�u�w�8��ԜY���F��F��*���r�#�;�u�9�}�������W������u�u�u�u�w�4�Wǿ�&����F�G�����u�u�u�u�w�}�W���	�֓�V ��[��*���2�i�u�%�4�3����J����9F�N��U���u�9�0�u�w�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������_��h�����u�;�u�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO�G�����_�u�u�u�w�}�W���Y���C9��E�����4�%�0�u�j�-�G�������[��N��U���u�u�u�u�2�9���s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����^��V�����'�2�4�&�0�}����
���l�N��D���3�8�-�4��1�(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���
�4�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��E�������9F�N��U���u�u�u�u�w�}�W���&����^��V�����'�2�i�u�'�>��������lV��N��U���u�u�u�u�w�}�����έ�l��h��*��u�=�;�_�w�}�W���Y���F�N��Uʥ�d�'�3�8�/�<�(���&����Z�G1�����8�-�4�
�;�f�W���Y���F�N��U���;�u�3�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*ۊ�0�
�4�
�%�:�����Ƽ�\��D@��X���u�%�d�'�1�0��������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��D���3�8�-�%�2�}�JϿ�&����G9��\��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�}�'�>��������lW������6�0�
��$�l����I�ƭ�WF��G1�����9�2�6�e�j�<�(��������F��*���&�
�:�<��}�W���&����^��V�����|�!�0�u�w�}�W���Y���F�N��*ۊ�0�
�4�
�%�:�K���&¹��U9��OUךU���u�u�u�u�w�}������ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�]�}�W��	�ԓ�V��S1��*���
�'�2�4�$�:�W�������K��N������'�:�
�'�+��������@��h����%�:�0�&�6�����Y����V��=N��U���u�3�}�%�4�6����Ӈ����T��H���d�|�!�0�]�}�W���Y���Z �V�����u�d�|�!�2�W�W���Y���F�N��G���'�:�
�%�!�9����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F�N��U���u�u�u�3��<�(���
����T��N�����0�|�!�0�]�}�W���Y���F�N�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��E�������9F�N��U���u�u�u�u�w�}�W���&����\��G1�����0�u�h�4��2��������]ǻN��U���u�u�u�u�w�}����Yۇ��@��U
��B���!�0�u�u�w�}�W���Y���F�N��U���
�0�<�1�6��������F��1�����
�%�#�1�]�}�W���Y���F�N�����<�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�G1��%���:�
�'�2�6�.��������@H�d��Uʥ�g��'�:��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h>�����%�0�u�h�6�����&����lV��N��U���u�u�0�&�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u����������E
��G�����_�u�u�u�w�}�W���Y���C9��g�����'�2�i�u���������F�N��U���u�0�1�<�l�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߠu�u�x�u����������C9��S1�����&�<�;�%�8�8����T�����h��*���4�4�
�9��/����
����C��T�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�N��R���=�;�u�u�w�}�W�������C9��CN��R��u�=�;�u�w�}�W���Y�����h��*���4�4�
�9��/���Y����\��h�����n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�f�3�8�e�t�W������F�N��U���u�u�u�u�w�-�B�������R9��h��*���2�i�u�%�4�3��������l�N��U���u�u�u�u�w�8����Q����Z��S
��M���=�;�_�u�w�}�W���Y���F�N�����'�3�7�!��-����	����[��h[�����0�4�4�
�;�f�W���Y���F�N��U���;�u�3�_�w�}�W���Y���F��SN��N�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƓF�C��*ߊ�0�
�0�4�'�8�W�������A	��D�X�ߊu�u�
�
�2�����	����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N�����'�3�7�!��/���Y����\��h��G��_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�;�!��<�(���
����T��N�����<�
�&�$���ށ�
������F��*���&�
�:�<��}�W���
����O�V ��]���6�;�!�9�0�>�F��	�ӓ�V ��R�����9�|�|�!�2�}�W���Y���F�N��U���
�
�0�
�2�<����Y����lS��R�����_�u�u�u�w�}�W���Y����Z ��=N��U���u�u�u�;�w�;�}���Y���V��^�U���0�1�%�:�2�.�}�ԜY�����[�����:�%�&�'�0�n�DϿ�
����C��R��U���u�u�<�
�>���������A��V�����2�
�'�6�m�-����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�l�^Ϫ����F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-��������`2��C\�����g�|�u�=�9�W�W���Y���F�N��Uʼ�
�<��'��2�(������� F������:�
�:�%�f�i����J����9F�N��U���u�u�u�9�>�}�_�������l
��^��U���%�&�2�6�2��#���Hʹ��^9��G�����_�u�u�u�w�}�W���Y���Z*��^1�����:�
�
�0��e�W������]��[��E�ߊu�u�u�u�w�}�W����ƥ�l�N��U���u�0�1�<�l�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�W���T�ƭ�@�������{�x�_�u�w�/����Yۇ��P
��=N��U���<�_�u�u�w�}����	������Y�����%�6�>�h�p�z�W������F�N��U���}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��C���Y����9F�N��U���u�u�u�g�e�/���O��� ��1��*��b�%�n�u�w�}�W���Y��� ��E��G��u�h��
�"�d�D���B���F�N��U���u�6�%�
�2��N��E�ƥ�^��Q��Lߊ�g�_�u�u�w�}�W���Y�ƥ�]��1����a�u�h�<�2��(ށ�����9��X����!�u�f�n�w�}�W���Y���F��D ��*���
�m�g�i�w�/�������� 9��X����!�u�f�n�w�}�W���Y���F��V ��*܊�0�
�l�e�k�}����&Ź��lW��1��N���u�u�u�u�w�}�WϬ�H����lT��N�U���
� �d�e��o�}���Y���F�N�����d�d�'�2�e�e�W������W��B1�Eӊ�d�_�u�u�w�}�W���Y�Ƹ�C9��1����m�u�h�!�'�l�C���&����l��=N��U���u�u�u�u�w�0�(�������
V��S�����d�3�
�c��o�}���Y���F�N�����d�
�0�
�n�i�K�������l ��Y����u�u�u�u�w�}�W�������9��P1�@���h�!�%�`��(�F��&����F�N��U���u�u�!�%�b�����@���F��G1�*���d�e�
�g�]�}�W���Y���F�C��Cي�0�
�l�g�k�}����J����
P��G_�U���u�u�u�u�w�}����Aǹ��T9��X��Hʡ�%�m�
� �f�o�(��s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�����Ƽ�\��D@��X���u�%�:�0�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�d�|�!�2�W�W���Y���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�~�)��ԜY���F�N��Uʇ�;�0�
�9��3��������A��^�U���;�0�
�;�����K����9��h_�D���n�u�u�u�w�}�W���Yӂ��V��h�����0�
�e�m�k�}��������A	��Q��B���%�n�u�u�w�}�W���Y����l_��S�����
�d�'�2�d�i�W��	����W��E	��*���3�
�g�d�'�f�W���Y���F�N��*���g�d�
�0��m�O��Y����_T��1��*��d�%�n�u�w�}�W���Y�����V��A���2�g�l�u�j�-�!���&ǹ��lW��1��N���u�u�u�u�w�}�Wϭ�����P��R	��E��i�u�0�
�:�o�(���H����CT��N��U���u�u�u�u�#�-�(���&����Z�C��*���d�b�
�g�]�}�W���Y���F�C��F݊�0�
�e�f�k�}����N����S��h����u�u�u�u�w�}�W�������D9��E��F��u�h� �1�%�1� �������^��UךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��ԶY���F��D��U���6�&�{�x�]�}�W���������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�P���Y����9F�N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�n�;���P�Ƹ�VǻN��U���u�u�u�u�8�1����6����A��R����� �9�&�'�0�o�E���Dӄ��_9��r�����0�!�'���,����&����W��UךU���u�u�u�u�w�}�$���*����l'��X�����9�0�l�
�2��O��E�ƪ�l'��O!��*���:� �0��;�8�N؁�����l��=N��U���u�u�u�u�w���������G��C��*���'�2�g�l�w�`��������V9��E�� ���b�
� �a�e�-�L���Y���F�N��U���
�m�'�2�e�m�W������9��h[�*��_�u�u�u�w�}�W���Y����9��P1�E���h�!�%�m�1��G݁�K���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϿ�
����C��R��U���u�u�%�:�2�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�d�|�#�8�}���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���g�3�8�g�~�t����s���F�N��U���6�
��������K�Г�lW��R	��E���i�u�!�e�c�h������ƹF�N��U���u�u�!�e�c�h��������A��^�U��9�
�
�a���(��s���F�N�����<�n�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�����Ƽ�\��D@��X���u�%�:�0�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�d�|�!�2�W�W���Y���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�l�|�w�5����Y���F�N��U���6�
�4�0��/��������9��P1�F���h�3�
�!��.�(�������V9��hZ�� ��b�%�n�u�w�}�W���Y��� ��T������'�6� �2�n�(܁�����T�
N��*����&�
�!�"�)����A�Փ�F9��1��N���u�u�u�u�w�}�Wϸ�&����R��d�����0�a�
�
�2��O��E�ƪ�l��t��*��� �!�'�
�b�i����Mʹ��l�N��U���u�u�u�3��)�4���&����P��R1�*ي�0�
�m�g�k�}�$���&����l5��B�����g�f�3�
�e��D�ԜY���F�N��Uʦ�9�!�%�
�2��O��E�ƿ�_9��G]�� ��d�%�n�u�w�}�W���Y�����T������'�6� �2�l�A�������F������4�0��'�4�(���O����
T��G]�U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K��D��ʥ�:�0�&�u�z�}�WϮ�����N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W��PӒ��]l�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�����P����[��N��U���u�u�u�u�1�����
����A��B��Fۊ�
�0�
�b�o�a�W���&����T��UךU���u�u�u�u�w�}�$���0����G9��1����m�u�h�2�'�;�(��&����F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W������]F��X�����x�u�u�%�8�8����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�d�~�)��ԜY���F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�f�3�8�f�t�^Ϫ����F�N��U���u�3�
�:�2�)����MĹ��T9�� _��Hʲ�%�3�
�g��l�}���Y���F�N��������!��9�F�������Q��S����� �f�`�%�l�}�W���Y���F������,� �
�1��m�(���&����Z�P�����l�
�g�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dךU���x�4�&�2�w�/����W���F�G�����}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�I�����_�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���!�0�_�u�w�}�W���Y���U5��z;�����
� �!�%�.�l�B�������F��������!��;�4����Kƹ��lR��h����u�u�u�u�w�3�W���s���F�R ����u�u�0�1�'�2����s���K�V�����'�6�&�{�z�W�W�������@F��G1���ߊu�u�0�<�]�}�W���Y���R��[�����u�;�u�%�4�6�J���^�Ƹ�VǻN��U���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o�(���&���F��R ךU���u�u�u�u�w�}�;���&����	��h_�*���
�e�a�i�w���������\��Z�� ��m�
�g�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dךU���x�4�&�2�w�/����W���F�G�����}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�I�����_�u�u�u�w�}�W���Q����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\ʺ�u�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��D���PӒ��]l�N��U���u�u�u�'�0�i�@��Y����U��]��G�ߊu�u�u�u�w�}�������F�N��ʼ�n�u�u�0�3�-����
��ƹF�N�����u�'�6�&�y�p�}���Y����V�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���^���G��=N��U���u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�E߁�
����F��SN�����:�1�3�
�a�n����Y����\��h��*���|�!�0�_�w�}�W���Y���F��G1�*���
�e�l�e�w�`����@����lT��1��]���_�u�u�8��n����J����O�
N����
� �g�l��l�F��Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�u�u�z�}����Ӗ��P��N����u�'�6�&�w�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����r�r�u�=�9�}�W���Y�����F�����;�!�9�2�4�l�JϿ�&���R�������!�9�2�6�f�`��������V��c1��Dӊ�&�
�m�|�w�5����Y���F�N��U���6�
�4�0��/��������l��C1����`�}�|�i�w���������G��C��*��
�4�!�3��k�G���Q����F�B,�����&�
�!� �#�/�(��&����l��h]�C��u�h� �
�$���������F��Z�����
� �g�m��l�F��Y����q9��h-�����'�6� �0�f�k����&���� V��\��I����6�
�4�2���������P��V�����c�e�%�}�~�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߊu�u�x�4�$�:�W�������K��N�����0�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��D���!�0�_�u�w�}�W���Y���N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l�� 1����|�|�!�0�]�}�W���Y���F�B"�����&�
�!� �#�/�(��&���� V��R�� ���!��&�
�#�(����&����U��^����u�u�u�u�w�}�W�������l%��R1����� �0�d�c�%�:�D��Y����9��h-�����'�6� �0�f�k����O�֓� ]ǻN��U���u�u�;�u�1�W�W���Y�Ʃ�WF��d��Uʰ�1�%�:�0�$�W�W���;����p��h=�� ���'�
�a�
�6�)����J����F��@ ��U���i�u�e�e�g�f�W������� 9��P1�C���f�1�"�!�w�t�K���I����V��^�E��e�e�e�e�g�m�G��I����V��^�E��e�e�e�e�g�m�U�ԶY���F��RN�����!�!�u�4������Y����[��C��U���=�;�{�x�]�}�W���7����^9��D��*���6�o�%�:�2�.�_���:����^J��G1��Yʴ�
�<�
�1��n�[ϻ�����W9��h\�F���|�u�u�7�0�3�W���Y����R��V��&���8�<�_�u�w�}�W���Y������d:��ۊ�&�
�u�k�]�}�W���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����%�&�2�7�3�l�E���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:��؊�&�
�n�u�w�}�W���Y�����Rd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�d�3�8�g�W�W���Y���F�N��ʼ�n�u�u�u�w�}�Wϩ��ƭ�l5��D�����d�h�u�u�w�}�W���Y�����y=�����h�4�
��$�n����K���F�N��Uʢ�0�u�%���)�(���&���l�N��U���u�u�u�4������E�ƭ�l5��D�����f�_�u�u�w�}�W�������C9��h��*���
�u�k�_�w�}�W���Y���F��h �����i�u�%���)�(���&��ƹF�N��U���=�;�4�
��.�B������FǻN��U���u�u�u�u�'��(���Y����C9��h��*���
�n�u�u�w�}�W�������R��c1��C���8�`�h�u�w�}�W���Y���F��G1��*���u�h�4�
��.�@�������F�N��U���"�0�u�%���؁�
����X�N��U���u�u�u�u�6��$������R��c1��M���8�b�_�u�w�}�W���Y������d:��Ҋ�&�
�u�k�]�}�W���Y���F�V��&���8�i�u�%���ց�
����9F�N��U���u�=�;�4��	��������[�=N��U���u�u�u�u�w�-�9���
�����d:�����3�8�l�_�w�}�W���Y�ƻ�V��G1��*���e�3�8�l�j�}�W���Y���F�N�����
�&�u�h�6��#���H¹��^9��d��U���u�u�u�"�2�}����&����l ��h_�H���u�u�u�u�w�}�W�������l ��R������&�d�
�$��F�ԜY���F�N�����%��
�!�e�;���Y���F�N��U���u�u�4�
��;���Y����g9��]�����g�_�u�u�w�}�W�������C9��h��F���8�d�u�k�]�}�W���Y���F�V��&���8�i�u�%���������� ]ǻN��U���u�u�=�;�6��#���Hǹ��^9��S����u�u�u�u�w�}�W���7����^F���&���!�`�3�8�f�f�W���Y���F��_������&�d�
�$��C��Y���F�N��U���u�%��
�$�}�JϿ�&����GW��Q��D��u�u�u�u�w�}� ���Y����g9��X�����`�h�u�u�w�}�W���Y�����y=�����h�4�
��$�l�(���&����F�N��U���"�0�u�%����������F�d��U���u�u�u�u�w�<�(������F��h=����
�&�
�b�]�}�W���Y���D����&���!�m�3�8�f�}�I�ԜY���F�N��Uʴ�
��3�8�k�}����&����l ��h_����u�u�u�u�w�5�Ͽ�&����GW��Q��D���k�_�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!�g�;���B���F�N��U���;�4�
��$�o�(���&���FǻN��U���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�3��������]��B1�Mي�g�h�4�
�8�.�(���&���F��R ךU���u�u�u�u�w�}�W���	����U��S�����
�!�g�3�:�o�L���Y���F�N��U���0�u�u�u�w�}�W���Y�����y=�����h�4�
��$�o�(���&����F�N��U���u�u�0�1�>�f�W���Y���F��_������&�g�
�$��G��Y���F�N��U���u�%��
�$�}�JϿ�&����GT��Q��D��u�u�u�u�w�}� ���Y����g9��\�����d�h�u�u�w�}�W���Y�����y=�����h�4�
��$�o�(���&����F�N��U���"�0�u�%����������F�d��U���u�u�u�u�w�<�(������F��h=�����3�8�e�_�w�}�W���Y�ƻ�V��C����u�_�u�u�w�}�W���Y�ƭ�l(��Q��I���������/���!����k>�=N��U���u�;�u�4�2�W�W����Ƽ�\��DUךU���g�g�3�
�g�j����Dӕ��l
��^�����'� �&�2�2�u��������EW��]�U���;�<�;�1�#�-�Cց�����9��G�U���u�u��
��<����&����l��S�����:�<�
�0�#�/�����ο�T��(��A���
�g�`�%�~�n�^��s���uT��h��D��
�f�i�u�w�}�W���?����T9��]�����}�8�
�f�1��E���	����[�I�����u�u�u�u�w�)���&����R��G\�U���u�u��
��<����&����l��S�����:�<�
�0�#�/�����ο�T��(��@���
�b�l�%�~�n�^��s���uT��h��D��
�f�i�u�w�}�W���?����A��W�U���;�}�8�
�d�;�(��@����O�I�\ʰ�&�u�u�u�w�}����Lƹ��lW��1��N���u��
� �n�n����Dӕ��l
��^�����'� �&�2�2�u��������EW��]�U���;�<�;�1�#�-����&����CW�d��Uʇ�;�0�
�9��3��������
U��N�U¡�%�
� �d�o��EϿ�Ӓ��lU��Q��@���%�|�_�u�w�<��������]��1��*��`�%�u�h��<��������]��1��*���g�f�
�f�6�9�%���¹��_9��R��*���g�b�
�g�l�}�Wό�����R
��X ��*؊�d�d�
� �e�i�(��E����R��h_��D���
�e�b�%�w�3�W����ד�_
��Y��G���
� �g�d��n�L���YӴ��T��V�����
�
�d�3��o�E���Y���F�N��'���0�
�9�
�9�.�E���&����l��@��Uº�
�:�1�f�>����Jʹ��V�
N��R���9�0�_�u�w�}�W���&����9��h\�A���n�u�u��9�8�(���&����lT��h_�����b�d�%�u�j�u����&¹��U��\�����;�u�4�2�f�<��������Z9��h_�L���|�_�u�u�6�:�F�������@9��^1��*��l�%�u�h�]�}�W���Y����VW��[�����3�
�c�d�'�}����Q����\��1�����c�`�%�}�~�`�P���Y����l�N��Uʦ�9�!�%�a�1��@���	��ƹF��V ��D���9�:�0�
��(�E��&���F��Z�����e�g�%�u�9�}����L����V��h�N���u��;�0��1�(���
����P��h�I����;�0�
�;�����H����F9��Y��Fʴ�1��;�0��1�(���
�ד�F9��]��G��u�u��;�2���������9��h_�D���u�h�w�w� �8�Wǳ�����F9��V��F��4�
�:�&��+�C��Y����D��d��Uʇ�;�0�
�9��8����&����S��G\��H���4�2�d�4�;�2����&����Q��G\�����%�6�;�!�;�l�F��Y����R��1�����'�&�g�<��(�E��&���FǻN��U���
�m�<�
�"�o�A܁�Kӑ��]F��E1����
�d�3�
�f�d����P���A�R��U���u�u�u�&�;�)��������V��UךU���4�2�d�4�;�'����K����F9��[��F��u�u�u�u�w�-�Nׁ�&����Q��G\�����}�'�6�;�n��(���H����CT�N��R��u�9�0�_�w�}�W�������CT��Q��B���%�n�u�u��3�ށ�����A	��1��*��`�%�u�h�u�� ���Yۋ��l0��h��*��e�h�4�
�8�.�(���M���V
��L�N���u��;�0��1�(�������lW��1��U��}�4�2�d�6�1����&¹��lW��1��U���u�%�6�;�#�1�F��B���4��P��#���3�
�c�l�'�}�Jϭ�����Z��R��¦�<�!�'�2�#�(�����Ρ�]9��Q��G���%�|�!�
�9�8��������V�I��U���
�a�3�
�a�h����H����\��XN�\���n�u�u��9�8�(���&����W��G\��Hʦ�1�9�2�6�!�>��������A��CF�����0�}�4�
������@���G	��Y�����;�<�;�1�p�z�QϪ�	����U��_�����d�d�1�"�#�}�^���P���F��Y	��*���
�;�&�d�1��F���	���D�������4�2�g��d�;�(��M����F��a1�����d�l�%�|�2�.�W��B���4��P�����:�0�
�
�f�;�(��H����[�N��U����;�0�
�;�����H����W��h����u�:�
�:�3�l�ށ�����9��^��H��r�u�9�0�]�}�W���Y����l ��^�*��_�u�u�4�0�o��������9��Q��C���%�u�h�_�w�}�W�������l��h�����
�c�d�%�w�5��������W_��^1��*��l�%�}�|�j�z�P������F�N�����
� �d�e��o�}���Y����VT��[�����3�
�c�d�'�}�J���[ӑ��]F��V ��G���d�3�
�c�n�-�W���&����lW��1��\ʰ�&�u�e�n�]�}�W������]��D��ʥ�:�0�&�u�z�}�WϿ�&����l��^	�����u�u�'�6�$�u����UӇ��@��T��*���&�g�
�&��o�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�f�1�0�E���PӒ��]FǻN��U���u�u�%�1�9�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʴ�
�1�0�4�$�:�W�������K��N�����1�0�4�&�0�����CӖ��P�������!�u�%�&�0�>����-����l ��h^��U���7�2�;�u�w�}�WϷ�Y�΢�GN��G1�����9�2�6�d�j�<�(������R�������!�9�2�6�f�`��������V��c1��D���8�e�|�u�?�3�}���Y���F�V�����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϿ�&����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��V
�����2�u�'�6�$�s�Z�ԜY�ƭ�l��S�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�e�����K���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�D�������O��_�����u�u�u�u�w�-���� ���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�'�4�,�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����u�:�;�:�`�t�}���Y����C��R���ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����f�1�"�!�w�n�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��\�����;�%�:�u�w�/����Q����G��N��E���3�4�%�4�6���������F��1�����-�4�
�9��3����Y����c��X
�����1�<�
�<�{�-�B�������R9��h��*���&�2�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��n�W��Qۖ��l��h�����
�9�
�;�$�:�JϿ�&����G9��P��E���'�}�
�
�2�4����&����Z��^	��U���6�;�!�9�0�>�G����μ�9��Q1�����
�9�
�;�$�:�JϿ�&����G9��P��E���'�}�
�
�2�����&����_��Y1����4�
�:�&��2����PӉ����D����4�
�:�&��2����P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��W�����;�%�:�0�$�}�Z���YӇ��@��U
��D���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�d�l�k�}��������_��N������3�8�c�3�*����P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��_�����;�%�:�0�$�}�Z���YӇ��@��U
��D���4�&�2�
�%�>�MϮ�������t=�����u�u�7�2�9�}�W���Y���F������7�1�d�d�k�}��������_��N������3�8�m�3�*����P��ƹF��Y
�����&�n�_�u�w�p�W���
����W��]����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��`�4�&�2��/���	����@��G1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�d�d�}�J���	����@��A_��U���%��
�&��}�������l�N��ʥ�:�0�&�_�]�}�W������T9��S1�A���&�<�;�%�8�8����T�����D�����d�a�
�&�>�3����Y�Ƽ�\��DF��*���3�8�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��k�D��Yۇ��P	��C1��D��h�4�
��1�0�EϺ�����O�=N��U���u�'�6�&�l�W�W���T�ƭ�l��h��*��d�4�&�2�w�/����W���F�V�����1�
�c�d�6�.���������T��]����
�&�|�w�}�������F�N��U���u�%�&�2�5�9�F��Y���R��X ��*���
�u�u�%������Y����G	�G�U���0�1�%�:�2�.�}�ԜY�����D�����d�`�u�&�>�3�������KǻN�����2�7�1�d�b���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����O���F��G1�����9�d�d�h�6��$�������\��XN�\�ߊu�u�;�u�%�>���s���K�V�����1�
�c�c�6�.��������@H�d��Uʴ�
�<�
�1��k�A���
����C��T�����&�}�%���.�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������F�F��*���&�
�#�
�w�}����&����F��@ ��U���n�u�u�0�3�-����
��ƓF�C�����2�7�1�d�n�<����Y����V��C�U���4�
�<�
�3��@ց�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������
F�F��*���&�
�#�
�w�}����&����
F��@ ��U���n�u�u�0�3�-����
��ƓF�C�����2�7�1�d�n�<����Y����V��C�U���4�
�<�
�3��Nց�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������
F�F��*���&�
�#�
�w�}����&����W��X����|�n�u�u�2�9��������9l�N�U���&�2�7�1�e�d�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����V��S�����:�&�
�#��}�W���:����^N��
�����d�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�o�BϿ�
����C��R��U���u�u�4�
�>�����Kƹ��@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9��N�U´�
�:�&�
�!��W���	����U��Z�����:�d�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�E������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��X�I���4�
�:�&��+�(���Y����`9��ZF�U���;�:�d�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���@Ӈ��Z��G�����u�x�u�u�6���������
9��D��*���6�o�%�:�2�.����*����l�N�����u�u�u�u�w�}�W�������T9��S1�L��u�4�
�:�$��ށ�Y�ƭ�l%��Q��D���:�;�:�d�~�f�W�������A	��D����u�x�u�%�$�:����J����@��YN�����&�u�x�u�w�<�(���&���� V��V�����'�6�o�%�8�8�ǿ�&����@�N�����;�u�u�u�w�}�W���YӇ��@��U
��F��i�u�4�
�8�.�(���&���R��d1����u�:�;�:�f�t�L���YӃ����T��N�ߠu�u�x�u�'�.����������^	�����0�&�u�x�w�}��������W9��1�����
�'�6�o�'�2��������l ��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����d�i�u�4��2����¹��F��h-�����d�u�:�;�8�l�^��Y����]��E����_�u�u�x�w�-�������� S��D��ʥ�:�0�&�u�z�}�WϿ�&����Q��]�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����f�`�i�u�6�����&����F�V��&���8�g�u�:�9�2�E���B����������n�_�u�u�z�}��������lU��V�����'�6�&�{�z�W�W���	����l��h]�����2�
�'�6�m�-����
ۇ��p5��D��U���7�2�;�u�w�}�W���Y�����D�����f�u�h�}�'��(���Q�ƨ�D��^��Hʴ�
�:�&�
�!��^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6���������F��D��U���6�&�{�x�]�}�W���
����W��\�����;�%�:�u�w�/����Q����`9��ZGךU���0�<�_�u�w�}�W���Y���R��^	�����l�u�h�}�'�>�����ד�[��G1��*���}�e�1�"�#�}�G���s���V��G�����_�_�u�u�z�<�(���&����V��V�����'�6�&�{�z�W�W���	����l��hZ�*���<�;�%�:�w�}����
�έ�l%��Q�����u�0�<�_�w�}�W���Y���F��h��*���
�e�u�h��-��������lW���6���&�}�b�1� �)�W��P���F��SN�����&�_�_�u�w�p��������W9�� N�����u�'�6�&�y�p�}���Y����Z��S
��D݊�&�<�;�%�8�}�W�������R��d1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�d�u�j�u��������EW��S�����
�&�}�g�3�*����K����F�R �����0�&�_�_�w�}�ZϿ�&����Q��]����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*��
�&�<�;�'�2�W�������@N��h-�����_�u�u�0�>�W�W���Y���F�N��*���
�1�
�f�w�`�_�������l
��h_��U����
�&�}�g�9� ���Y���l�N��ʥ�:�0�&�_�]�}�W������T9��S1�U���<�;�%�:�2�.�W��Y����C9��P1�����
�&�<�;�'�2�W�������@N��h�����4�
�<�
�$�,�$���¹��^9����*���
�9�=�
�'�+��ԜY�Ʈ�T��N��U���u�u�u�u�6���������Z�F��*���&�
�:�<��}�W���&����R
��V1��*���|�4�1�;�#�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��Y
�����:�&�
�:�>��W���	����A�G�U���0�1�%�:�2�.�}�ԜY�����D�����c�u�&�<�9�-����
���9F������7�1�c�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
�0�
�6��������F��P��U���u�u�u�u�w�}��������W9��R��]���}�}�%�6�9�)���������D�����
��&�d�1�0�G�������C9��Y�����6�e�h�4��)����PӇ��N��h�����:�<�
�u�w��(���&����R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�b�u�&�>�3�������KǻN�����2�7�1�b��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�0�>�9������ƹF��R	�����u�u�u�u�w�}�W���
����W��N�U»�!�}�4�
�8�.�(�������F��h��*���$��
�!��.�(������R��X ��*���<�
�u�u�'�.����P�ƭ�WF��G1�����9�2�6�d�j�-�E�������R��[
��N���u�0�1�%�8�8��Զs���K��G1�����1�m�u�&�>�3�������KǻN�����2�7�1�m��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�0��8����&����9F����ߊu�u�u�u�w�}�W���	����l��hV�I���;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`��������V��V�����n�u�u�0�3�-����
��ƓF�C�����2�6�0�
��.�F߁�
����R��P �����&�{�x�_�w�}��������B9��h��E���8�l�4�&�0�����CӖ��P�������7�1�d�l�]�}�W������F�N��U´�
�<�
�1��j�^Ϫ���ƹF�N��U���%�&�2�6�2��#���Hù��^9��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��h��*���h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���&�2�6�0��	���&����V��D��ʥ�:�0�&�u�z�}�WϿ�&����P��h=����
�&�
�e�6�.���������T��]���&�2�7�1�c�d�}���Y����]l�N��Uʼ�u�4�
�<��9�(��PӒ��]FǻN��U���u�u�%�&�0�>����-����9��Z1�U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}��������B9��h��D���8�d�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�>����-����9��Z1�U���<�;�%�:�2�.�W��Y����C9��P1������&�d�
�$��F���
����C��T�����&�}�%�&�0�?���@���F��P��U���u�u�<�u�6���������
O��_�����u�u�u�u�w�-��������`2��C_�����d�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����Z��D��&���!�g�3�8�f�}�JϿ�&����G9��P��E�ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w�-��������`2��C_�����d�u�&�<�9�-����
���9F������6�0�
��$�l�(���&�ԓ�@��Y1�����u�'�6�&��-��������_�N�����;�u�u�u�w�4�Wǿ�&����Q��^�U���;�_�u�u�w�}�W���	����l��F1��*���f�3�8�d�w�`��������_	��T1����u�u�u�9�2�W�W���Y���F��h��*���$��
�!�d�;���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��F1��*���a�3�8�d�w�.����	����@�CךU���%�&�2�6�2��#���Hǹ��^9��h�����%�:�u�u�%�>����	����l��h_�\���u�7�2�;�w�}�W�������C9��P1����b�u�=�;�]�}�W���Y���R��^	������
�!�a�1�0�F���DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����<�
�&�$���������� F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��^	������
�!�`�1�0�F���
������T��[���_�u�u�%�$�:����&����GW��Q��Dފ�&�<�;�%�8�}�W�������R��^	�����g�|�u�u�5�:����Y����������7�1�g�`�w�5��ԜY���F�N��*���
�&�$���)�B�������[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����l ��h_�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���
�&�$���)�A�������R��P �����&�{�x�_�w�}��������B9��h��C���8�d�
�&�>�3����Y�Ƽ�\��DF��*���
�1�
�c�~�}�Wϼ���ƹF�N�����%�&�2�7�3�o�D������F�N��U���4�
�<�
�$�,�$����Г�@��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����
����g9��X�����`�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�<�
�$�,�$����ѓ�@��N�����u�'�6�&�y�p�}���Y����Z��D��&���!�b�3�8�f���������PF��G�����4�
�<�
�3��O���Y����V��=N��U���u�3�}�%�$�:����K���G��d��U���u�u�u�4��4�(�������@��h��*��i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϿ�&����P��h=����
�&�
�c�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��h��*��4�&�2�u�%�>���T���F��h��*���$��
�!�o�;���&����T��E��Oʥ�:�0�&�4��4�(���&����9F����ߊu�u�u�u�1�u��������lR��N�����u�u�u�u�w�}��������V��c1��DҊ�&�
�b�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�d�
�$��@��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��Dӊ�&�
�m�4�$�:�W�������K��N�����<�
�&�$����������9��D��*���6�o�%�:�2�.��������W9��GךU���0�<�_�u�w�}�W���Q����Z��S
��E���!�0�u�u�w�}�W���YӇ��@��T��*���&�d�
�&��e�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�l�(���&���F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�d�3�8�g�<����Y����V��C�U���4�
�<�
�$�,�$���¹��^9��V�����'�6�o�%�8�8�ǿ�&����Q��W��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��F���!�0�u�u�w�}�W���YӇ��@��T��*���&�d�3�8�g�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����0�
��&�f�;���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϿ�&����P��h=����
�&�
�l�6�.��������@H�d��Uʴ�
�<�
�&�&��(���I����lW��V�����'�6�o�%�8�8�ǿ�&����Q��_����u�0�<�_�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y����C9��P1������&�g�
�$��N��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�E߁�
����Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�g�
�$��GϿ�
����C��R��U���u�u�4�
�>�����*����W��D��E���&�2�
�'�4�g��������C9��P1����g�_�u�u�2�4�}���Y���Z �V�����1�
�l�|�#�8�W���Y���F������6�0�
��$�o�(���&���F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�&�2�4�8�(���
����U��^��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�o�(���&����@��YN�����&�u�x�u�w�<�(���&����l5��D�*���
�d�4�&�0�����CӖ��P�������7�1�f�`�]�}�W������F�N��U´�
�<�
�1��n�^Ϫ���ƹF�N��U���%�&�2�6�2��#���K����^9��R�����:�&�
�:�>��L���Y�����RNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���%�&�2�6�2��#���K����^9�������%�:�0�&�w�p�W�������T9��R��!���g�
�&�
�e�<����&����\��E�����%�&�2�7�3�i�@�ԜY�Ʈ�T��N��U���<�u�4�
�>�����H����[��=N��U���u�u�u�%�$�:����&����GT��Q��G���h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���
����@��d:�����3�8�g�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GT��D��U���<�;�%�:�2�.�W��Y����C9��P1������&�g�3�:�l��������\������}�%�&�2�5�9�F��P�����^ ךU���u�u�3�}�'�.��������O��_�����u�u�u�u�w�-��������`2��C\�����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GU��D��U���<�;�%�:�2�.�W��Y����C9��P1������&�f�3�:�o��������\������}�%�&�2�5�9�F��P�����^ ךU���u�u�3�}�'�.�������� O��_�����u�u�u�u�w�-��������`2��C]�����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GR��D��U���<�;�%�:�2�.�W��Y����C9��P1������&�a�3�:�n��������\������}�%�&�2�5�9�F��P�����^ ךU���u�u�3�}�'�.��������O��_�����u�u�u�u�w�-��������`2��CZ�����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GS��D��U���<�;�%�:�2�.�W��Y����C9��P1������&�`�3�:�i��������\������}�%�&�2�5�9�F��P�����^ ךU���u�u�3�}�'�.��������
O��_�����u�u�u�u�w�-��������`2��C[�����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GP��D��U���<�;�%�:�2�.�W��Y����C9��P1������&�c�3�:�h��������\������}�%�&�2�5�9�F��P�����^ ךU���u�u�3�}�'�.��������O��_�����u�u�u�u�w�-��������`2��CX�����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�%�$�:����&����GQ��D��U���<�;�%�:�2�.�W��Y����C9��P1������&�b�3�:�k��������\������}�%�&�2�5�9�F��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��h��*���h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W���
����@��d:��݊�&�
�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�>����-����l ��hY�����;�%�:�0�$�}�Z���YӇ��@��T��*���&�m�3�8�`�<����&����\��E�����%�&�2�7�3�l�O�ԜY�Ʈ�T��N��U���<�u�4�
�>�����I����[��=N��U���u�u�u�%�$�:����&����G^��D��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}��������B9��h��*���
�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
�ߓ�@�������%�:�0�&�w�p�W�������T9��R��!���l�3�8�m�6�.���������T��]���&�2�7�1�f�l�}���Y����]l�N��Uʼ�u�4�
�<��9�(��PӒ��]FǻN��U���u�u�%�&�0�>����-����l ��hV��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��CW�����u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǻN�����-���!��8����6����F��D1��*���
�g�i�u�#�-�C݁�����l��V �����a�
� �a�d�-�^�ԜY�Ʈ�^��R_�� ��e�
�g�i�w�(��������l��h��G��
�g�:�u��j��������ZU��h ��*���g�l�
�g�l�}�Wϼ�����l ��]�*��i�u� �1�%�1� �������U��h����
�b�1�8�%�<�(�������lT��1��\�ߊu�u�'�0�0��(��L����l ��]�*��i�u�%�l��8��������A��^�U���u�;�0�3�8��(���&���� ^��G\����u�'�0�2���(���&���� U��G\��H���
�b�1�8�%�<�(�������9����U���0�3�:�
�8����KĹ��]ǻN�� ���
�g�l�4�3�8����DӒ��l_��Q��C���%�}�u�u�w�2����I��ƓF�C�� ���
�g�l�4�3�8����
������T��[���_�u�u� ���E�������@��V�����'�6�o�%�8�8�ǿ�&����P��h=����
�&�
�c�w�-��������`2��C_�����d�y�4�
�>�����*����^��D��B�ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�6�����
����g9��W�����m�|�!�0�w�}�W���Y�����h^��G���4�1�0�&�w�`��������_��h\��U���u�:�;�:�g�f�W���Y����_��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�b�~�)����Y���F�N�� ���
�g�l�4�3�8����DӇ��P	��C1��Cފ�}�u�u�u�8�3���B���F������}�%�6�;�#�1����H����C9��P1������&�d�
�$��A�������9F�N��U���u� �
�
�e�d��������[��G1�����9�c�
�}�w�}�W������]ǻN��U���9�0�_�u�w�}�W���Y����9��W�����&�d�i�u���}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��Q1��D��
�0�u�&�>�3�������KǻN�� ���
�g�l�6�g�<����&����\��E�����%�6�y�4��4�(�������@��h��*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C\�����d�|�|�!�2�}�W���Y���F��B��*��l�6�e�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����F ��h_�L���e�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���7�3�e�d�c�����
������T��[���_�u�u� ���E����ד�@��Y1�����u�'�6�&��-�������T9��R��!���d�
�&�
�a�}��������B9��h��L���8�d�y�4��4�(�������@��h��*��_�u�u�0�>�W�W���Y�ƥ�N������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�c�|�:�w�u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�Fց�
����O��EN�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�~�}����s���F�N�����e�d�a�
�2�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�U��E��a�
�0�u�j�<�(���
����T��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u� ���E����ƭ�@�������{�x�_�u�w�(�(߁�K�ߓ�9��D��*���6�o�%�:�2�.��������V9��E�� ���d�l�'�2�d�i�[Ͽ�&����P��h=����
�&�
�c�w���������G��C��*��
�0�
�e�f�}��������B9��h��L���8�d�y�4��4�(�������@��h��*��u��6�
�6�8�$�������lW��h��G��
�f�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�m�~�)����Y���F�N�� ���
�g�l�1�w�`��������V9��E�� ���d�l�'�2�d�i�L���Y�����^��]���6�;�!�9�0�>�F������T9��R��!���d�
�&�
�`�t����Y���F�N��U���
�
�g�l�3�}�Jϫ�&����R��d�����0�d�c�'�0�n�B��Y���F��[��U���%�6�;�!�;�:���DӇ��@��T��*���&�d�
�&��k�^Ϫ���ƹF�N��U��� �
�
�g�n�9�W������l%��R1����� �0�d�f�1��A���	��ƹF�N�����_�u�u�u�w�}�W���&ù��_��N�Uȍ�������/���!����k>��o6��-��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�?����H����D��V�����'�6�&�{�z�W�W�������T��h��*���<�;�%�:�w�}����
�έ�l�������6�0�
��$�l�(���&���R��^	������
�!�l�1�0�F������T9��R��!���d�
�&�
�`�W�W�������F�N�����}�}�%�6�9�)���������T�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��A������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���u�'�}�4��2��������F�V�����;�u�4�
�8�.�(�������F��h��*���$��
�!�o�;���P���G��d��U���u�u�u�7�1�m�F��&����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�7�3�e�f�i�(���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}����&¹��l ��^�*��i�u�!�%��(�E��&����]��R����
� �d�f��o�L���YӅ��A��h�� ��g�
�g�i�w�)����&����l��V �����!�%�`�3��i�C���P���F��V�����
� �a�e�'�}�Jϸ�&����g��C1�����9�
�g�
�2��O��s���W9��D��*���a�b�%�u�j�/���N���F��[�����'�&�d�3��o�A���Y���F�N��'���0�
�9�
�9�.�E���&����W��G]�����}�4�'�
��l����I�ѓ�N��S��D���0�&�u�u�w�}�Wό�����R
��M�����<�
� �g�e��D�ԜY�ƨ�_��S1�����3�
�b�f�'�}�J�ԜY���F��Y	��*���
�;�&�g�>�;�(��@����D��F�����d�<�3�
�b�l����P���A�R��U���u�u�u��9�8�(���&����@9��^1��*��`�%�n�u�w�8��������lT��1��U��w�w�"�0�w�4�(���?����\	��D1����f�h�4�
�8�.�(���&����_��^�����u�-�
�8���(���H����CR�
N�����
�
� �d�d��F��Y����G	�G�U���0�%�!�%��;�(��&���F��R	��*���l�f�%�}�e�9� ���Y���9F���4����!��&�;�)�(�������G	��B1�D���u�h�3�
��%��������G��V��*���g�3�
�c��n�}���Y����q5��B����� �0��9�2�d�(݁�����l��S��U���u�u�'�2�c�j� ���Yہ��l ��[�����|�h�r�r�w�1��ԜY���F��h/�����
�7�:� �2�����@Ĺ��lS��h����u�����)�6�������e��R1�*���`�e�%�u�j�;�(�������r��[��*��� �
�b�;�1��Bہ�K���F��h/�����
�7�:� �2�����@Ĺ��U��Z��G��u�3�
�!��.�(�������V9��h�����3�
�d�
�f�%�Ͽ�&����G9��\��E��e�e�n�u�w�;�(���:����`��T����
� �`�l�'�}�J�ԜY���F��h��6���
�!� �!�%��F�������Q��@��U²�%�3�
�a��o�G���Y�����RNךU���u�u��6��<��������A��1��*��
�d�_�u�w���������G��C��*���!�
�;�
�"�h�D���Y����`9��h-�����'�6� �0�e����@����9F������4�0��'�4�(���&ǹ��lQ��h�I���u�u�u�u�%�:�C��������h��F���
�l�
�g�g�}�W��PӃ��VFǻN��U����6�
�4�2���������9��Q��B؊�f�_�u�u��>�(�������F��E��D���3�
�g�
�d�a�W���Y��� ��T������'�6� �2�j�(���&������YN�����3�
�b�
�e�m�W���H����_��=N��U���u��6�
�6�8�$�������lU��Q��E؊�f�_�u�u��>�(�������F��E��D���3�
�a�
�d�a�W���Y��� ��T������'�6� �2�j�(���&������YN�����8�g�3�
�d��E��Y���O��[�����u�u�u��4�����*����G��h]��C���
�g�
�f�]�}�W�������@��C�����
�d�m�3��j�(��E��ƹF�N��&���
�4�0��%�>����J¹��A��Y�U���;�}�0�
�:�j����OŹ��V�
N��R���9�0�_�u�w�}�W�������@��C�����
�d�b�3��i�(��s���U5��C1�����!� �!�'��l����I����Z�=N��U���u��6�
�6�8�$�������lU��1����b�u�=�;��0�(ف�����l��G��U��|�0�&�u�w�}�W�������`��C1�����!�
�4� ��j����K����9F������4�0��'�4�(���&¹��l^��h�I���u�u�u�u�%�:�C��������h��G���
�f�
�g�g�}�W��PӃ��VFǻN��U����6�
�4�2���������9��hV�*��_�u�u��4�����*����G��h]��G���
�b�
�f�k�}�W���Y����`9��d�����&�9�!�
�6�(�(�������W��@��U¦�9�!�%�
�"�j�A���Q���A��N�����u�u�u�u�1�����
����A��B��FҊ�
� �m�f�'�f�W�������l%��R1����� �0�f�
��(�O���	���l�N��Uʳ�
��-� ��?��������F�� 1����d�u�=�;��8�(���J����_��G\��\��r�r�u�9�2�W�W���Y�ƪ�l��t��*��� �!�'�
�o�o����N¹��l�N��*����&�
�!�"�)����A����S��G]��H�ߊu�u�u�u���$�������\
��R1�����l�
�0�
�o�o� ���Yۏ��C9��hX�*��e�u�u�d�~�8����Y���F��R	��@��u�u�3�
�#���������F��[��*���m�l�%�u�j�W�W���Y�ƪ�l��t��*��� �!�'�
�e�/���@�ƻ�V�D�����
� �b�d�'�u�^��^���V
��d��U���u�&�9�!�'����K����9F������4�0��'�4�(���&¹��l^��h�I���u�u�u�u�%�:�C��������h��G���
�f�
�g�g�}�W��PӃ��VFǻN��U�������#���������_��Y�����m�g�_�u�w���������G��C��*���g�3�
�d��n�K���Y���F��R	��@���=�;�}�0��0�@���&����CT�N��R��u�9�0�_�w�}�W���*����p��h=�� ���'�
�g�d�1��Gځ�J���F��h��6���
�!� �!�%��E�������9��R�����u�u�u�0��h�W����ο�_9��G]�� ��d�%�}�|�j�z�P������F�N�����!��&�
�#�(����&�ԓ�l ��_����u�u�3�
�#���������F��\�� ��m�%�u�h�]�}�W���Y����S��@��U¡�%�c�3�
�n��E��Y���O��[�����u�u�u��4�����*����G��hY�����g�l�n�u�w�;�(���:����`��T�����
�:�<�!�1��F؁�H���A��[����u��6�
�6�8�$�������lQ��Q��B؊�d�i�u��4�����*����G��hY�����3�
�c�
�e�W�W���*����p��h=�� ���'�
�g�;�0�;�(��&���F��d1��*���0��'�6�"�8�@݁�����l ��X�����:�u�%�6�9�)���&����V��UךU����6�
�4�2���������9��h��*���a�f�%�u�j�;�(���:����`��T����
�
�0�
�`�e�}���Y����~3��N!��*���!�%�,�d�b�;�(��&���F��h��1���!��1�d�n�/���A��ƹF��d1�� ����!��9�>�1�(��&����^��N�U���;�1�
�0�:�i�@�������]ǑN��X���'�
� �f�b�>�W�������A	��D�X�ߊu�u�'�
�"�n�B���&����T��E��Oʥ�:�0�&�4��8�W���
����@��d:�����3�8�d�y�6�����
����g9��]�����g�u�%�&�0�>����-����9��Z1�\���u�7�2�;�w�}�W��������T�����2�6�d�h�6��������R��X ��*���<�
�u�u�'�.��������l��1����|�:�u�4��2��������F�V�����&�$��
�#�n����H����AF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�e�|�|�#�8�W���Y���F�	��*���f�`�6�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���T��Q��Lߊ�0�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]ǑN�����3�
�l�
�g�a�W�������@��C�����
�d�a�'�0�o�D��Y����A��B1�@���u�h�3�
�#���������F��\��*���
�m�g�_�w�}�Z�������lU��h�����2�u�'�6�$�s�Z�ԜY�ƫ�C9��h]�*���4�&�2�
�%�>�MϮ�������T����<�
�&�$����������J��G1�����0�
��&�f�����K�ƭ�l��h�����
�!�d�3�:�l�^���Yӄ��ZǻN��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�4�
�8�.�(�������F��h��*���$��
�!�e�;���PӉ����T�����2�6�d�h�6�����
����g9��]�����g�u�'�}�'�>��������lW������6�0�
��$�l�(���&���O��_�����u�u�u�u�w�/�(���J�ߓ�VF������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�2�%�1��Nց����R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}��������
9��R�����!��&�
�#�(����&�ӓ�l��h\�B�ߊu�u�'�
�"�n�N���Y����`9��h-�����'�6� �0�d��(���&����lǻN��Xʲ�%�3�
�e��m�����Ƽ�\��D@��X���u�2�%�3��m�(�������]9��X��U���6�&�}�%�$�:����&����G^��D��Yʴ�
�<�
�&�&��(���M����lW�������,� �
�d��8�(��@�ƪ�l��s�����1�d�c�'�0�o�@���Y����V��=N��U���u�3�}�4��2��������F�V�����&�$��
�#�i����H���G��d��U���u�u�u�2�'�;�(��&���F��h��1���!��1�d�a�/���N��ƹF�N�����u�}�%�6�9�)���������D�����
��&�m�1�0�@�������9F�N��U���u�'�
� �c�n����DӀ��K"��N!��*��
�0�
�b�n�W�W���Y�Ʃ�@�N��U���u�u�2�%�1��G܁�I���>��o6��-���������/���!����]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�'�
� �c�n����
������T��[���_�u�u�'��(�C���	¹��@��h����%�:�0�&�6�����
����g9��1����u�%�&�2�4�8�(���
����U��]����:�0�!�'��i�(���&����l�N�����u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���Hǹ��^9��G�����_�u�u�u�w�}�W���&����U��N�U���;�1�
�0�:�i�@�������]ǻN��U���9�<�u�}�'�>��������lW������6�0�
��$�e����N����[��=N��U���u�u�u�'��(�C���	�����T�����f�
��f��m�}���Y���V
��d��U���u�u�u�2�'�;�(��&���F��o6��-���������/���!����k>�=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�'�
�"�i�E���Y����T��E�����x�_�u�u�%����K����R��P �����o�%�:�0�$�<�(���&����l5��D�����e�u�%�6�{�<�(���&����U�������6�0�
��$�j����O�ƭ�l��h�����
�!�
�&��q��������V��c1��F���8�g�u�%�$�:����&����GR��D��Yʴ�
�<�
�&�&��(���&����J��G1�����0�
��&�a�;���s���Q��Yd��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�}�6�����&����P9��
N��*���
�&�$���)�(���&����]��X�����2�7�1�d�e�t��������]��[����h�4�
�<��.����&����U��G�����%�6�;�!�;�:���DӇ��@��T��*���&�g�3�8�f�}����	����@��X	��*���u�%�&�2�4�8�(���
�Փ�@��N��U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�2�Wǿ�&����G9��P��D��4�
�<�
�$�,�$���ƹ��^9����]���6�;�!�9�0�>�F������T9��R��!���c�3�8�`�~�t����Y���F�N��U���
� �a�g�4�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�P�����d�
�0�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���2�%�3�
�f��G��Y����A��V�����
�<�n�u�w�:����&����CW�
N��D���3�8�-�<��4�L�ԜY�����h��A���6�u�&�<�9�-����
���9F�	��*���a�m�6�
�$�4��������C��R�����<�
�&�$���ށ�
������T����<�
�1�
�d�q��������V��c1��B���8�c�u�%�$�:����&����GT��D��Yʴ�
�<�
�&�&��(���&����J��G1�����0�
��&�c�;���Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�����`�_�u�u�2�4�}���Y���Z �F��*���&�
�:�<��}�W�������]�F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�3�ǿ�&����Q��]�\ʺ�u�4�
�:�$�����&���R��^	������
�!�
�$��^ϱ�Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���}�%�6�;�#�1����H����C9��P1������&�f�3�:�o�W���Q����\��h�����u�u�%�&�0�>����-����l ��h]�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t��������]��[����h�4�
�<��.����&����U��G��\ʡ�0�u�u�u�w�}�W�������F9��1��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}��������l��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԜY�ƫ�C9��hZ�*��i�u�
�
�2���������T]ǻN����� �a�m�%�w�`��������R��Y1���ߠu�u�x�u�%����M����R��P �����&�{�x�_�w�}��������l��V�����'�6�o�%�8�8�ǿ�&���R��^	������
�!�g�1�0�F������T9��R��!���d�
�&�
�e�W�W�������F�N�����}�4�
�:�$�����&���R��RG�����}�%�6�;�#�1����H����C9��P1������&�d�
�$��F����έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���|�u�=�;�]�}�W���Y���T��Q��Gފ�0�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������F9��1��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƹF��E�� ��a�%�u�h�$�9��������G	��E�����;�<�;�1�'�o�'�������l��B�\��_�u�u�x�0�-����J����P	�������%�:�0�&�w�p�W�������F9��1�����
�&�<�;�'�2�W�������@N��h��*���$��
�!��.�(������T9��R��!���d�
�&�
�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�e�3�:�d�^Ϫ���ƹF�N��U���'�
� �a�d�2����Y����C9��Y�����f�_�u�u�w�}����Y�έ�l��D�����
�u�u�%�$�:����&����G_��D��\���=�;�_�u�w�}�W���Y����U��]�����0�i�u�%�4�3����L����F�N�����u�u�u�u�w�}�WϹ�	����U��X�����h�w���u�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����U��]��E��u��6�
�6�8�$�������lU��1����b�n�u�u�0�-����J����Z�V�����
�#�g�e�]�}�W��Y����U��V�����0�4�&�2�w�/����W���F�P�����f�
�%�:�2�<����&����\��E�����%�&�2�6�2��#���@����l^�V�����&�$��
�#�m����@���F��P��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�F߁�
����F��R ��U���u�u�u�u�0�-����J˹��P	��R�����:�&�
�#��f�W���Y����_��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�m�|�#�8�W���Y���F�	��*���a�m�:�6�3�}�JϿ�&����G9��1����u�u�u�9�2�W�W���Y���F��G1��*��
�%�:�0�k�}�/���!��ƹF�N�����3�u�u�u�2�9��������9F�	��*���a�m�%�u�j�/���N���F��G1��*��
�d�i�u�'�>��������]ǑN��X���'�
� �a�`�-�W�������A	��D�X�ߊu�u�'�
�"�i�@���&����T��E��Oʥ�:�0�&�4��4�(�������@��Q��M���8�
�
� �b�o�������l��h\�G���%�&�2�6�2��#���Hù��^9��=N��U���<�_�u�u�w�}��������]��[����h�4�
�<��.����&����l ��hW��U���;�_�u�u�w�}�W�������lR��h�I���8�
�
�0��e�E�ԜY���F��D��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}����s���F�N�����3�
�a�
�g�a�W���&˹��lS��h����u�u�u�9�2�W�W���Y���F��G1��*��
�e�i�u��f�W���Y����]��QU��U���0�1�%�:�2�.�}���YӁ��l ��Z�����h�}�'�
�"�i�@���Y����T��Q��Fي�g�n�_�u�w�p��������9�������%�:�0�&�w�p�W�������F9��1��*���<�;�%�:�w�}����
�έ�l��h�����
�!�
�&��q����H˹��lS��h�U���
�m�'�2�e�m�[Ͽ�&����P��h=����
�&�
�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�e�3�8�n�t����Y���F�N��U���
� �a�g�'�}�JϪ�	����A��V�N���u�u�u�0�$�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���ʹ��^9��N�����u�u�u�u�w�}��������9��R�����d�
� �`�`�-�L���Y�����RNךU���u�u�u�u�%����K����[�oL�U���u�u�0�1�>�f�}���Y����C��R�����u�2�%�3��h�(��E����A��B1�G���u�;�u�'��(�C���	����F�^"�����'��:�
�n����Aʹ��Z�D�����6�#�6�:��3����ۏ��_��X�����&�'�2�f�d�}�W���������T�����g�d�|�_�w�}����&����
S��N�U��u�=�;�}�>�3�Ǫ�	����U��[��A���u�<�;�1�6�����&����lV������w�_�u�u�4�-�(���H����CT�
N��Wʢ�0�u�!�%�f�o����A�Г�F�V�����
�#�
�|�2�.�W��B�����G]�� ��a�
�g�i�w�l�W����ο�T����*��
� �d�f��i�W���������T�����d�
�|�u�;�8�U���s���Z��1��*��c�%�u�h�u�� ���Yے��lP��Q��G���%�u�u�%�4�3����N���V
��L�N���u�<�8�
�"�k�D���Y���D��_��]���
�g�3�
�a��D������]��[��E���9�0�w�w�]�}�W���	����l �� [�����h�}�6�%�1��@܁�KӞ����T�����d�d�n�u�w�4����&¹��lW��1��U��1�4�&�2�����I����9F������3�
�f�
�f�a�W���
����l ��\����u�u�<�;�0�l����I�ߓ� F������d�3�
�e�f�-�_������\F��UךU����d�3�
�g�e����DӒ��lQ��Q��E���%�}�u�u�w�2����I��ƹF��s1��*���f�%�u�h�#�-�C߁�����9��_��U���:�;�:�e�l�W�W���Tӊ��9��1��E���1�0�&�u�$�4�Ϯ�����F�=N��U���e�a�`�0�g�<����
ù��@��h����%�:�0�&�6�����
����g9��^�����l�u�%�&�0�>����-����9��Z1�\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u�'�.��������l��1����|�u�=�;�]�}�W���Y���_��hZ�*���
�1�'�&�g�a�W�������l
��1�G���d�1�"�!�w�t�}���Y���V
��QN�����:�&�
�:�>��W���	����l��F1��*���e�3�8�d�~�}����s���F�N�����
�a�
�
��9����I���R��X ��*���a�e�g�x�f�9� ���Y����F�N�����u�u�u�u�w�}�Wϲ�&ù��9��1�����&�u�h�w��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY���
��1�@���e�4�1�0�$�}����Ӗ��P��N����u�!�e�a�b�8�G�������9��D��*���6�o�%�:�2�.����@����T9��W����<�
�&�$����������J��G1�����0�
��&�e�����I���F��P��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�Eށ�
����O��_�����u�u�u�u�w�)�G��L����l��E��D��u�8�
�f�%�:�D��Q���F��@ ��U���_�u�u�u�w�1����Q����\��h�����u�u�%�&�0�>����-����9��Z1�\���=�;�_�u�w�}�W���Y����lR��h��*���'�&�d�i�w�-��������9��N�Dʱ�"�!�u�|�]�}�W���Y����l�N��U���u�9�
�
�c��(߁�����@W�
N��-��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�1�(߁�Mƹ��9��N�����u�'�6�&�y�p�}���Y����lR��h��*���
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	���&����_�V�����&�$��
�#�o����K��ƹF��R	�����u�u�u�3��u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������
O�X��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�d�~�t����Y���F�N��U���e�a�`�0�g�>�G��Y����\��h�����n�u�u�u�w�8����Y���F�N�����a�`�0�e�4�m�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�1�(߁�Mƹ��9��N�����u�'�6�&�y�p�}���Y����lR��h��*���
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	���&����W�V�����&�$��
�#�l����K��ƹF��R	�����u�u�u�3��u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O�X��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�e�~�t����Y���F�N��U���e�a�`�0�g�>�F��Y����\��h�����n�u�u�u�w�8����Y���F�N�����a�`�0�e�4�l�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�u�u�9���Cځ�&ù��Z�B"��8���g��!�&�1��@���	��ƓF�C�����a�`�0�e� �l�����Ƽ�\��D@��X���u�9�
�
�c��(߁�¹��@��h����%�:�0�&�6�����	����l��F1��*���d�3�8�g�~�}�Wϼ���ƹF�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�d�3�:�o�^���Y����l�N��U���u�9�
�
�c��(߁������T�����2�6�d�_�w�}�W������F�N��U���9�
�
�a���(���Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z����֓�S��h_�����&�e�4�&�0�}����
���l�N��*ڊ�a�
�
�
�3�/��������]9��X��U���6�&�}�%�$�:����&����GT��Q��D���4�
�<�
�$�,�$����ԓ�@��GךU���0�<�_�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�>�����*����T��D��D���!�0�u�u�w�}�W���Yӊ��9��1��D���1�0�&�u�j�<�(���
����R��\��U���:�;�:�e�l�}�W���YӃ��Z ������!�9�2�6�f�`��������V��c1��Gڊ�&�
�l�|�#�8�W���Y���F���E��`�0�d�4�3�8����DӇ��P	��C1��Cފ�}�u�u�u�8�3���B���F����ߊu�u�u�u�w�}����M�ӓ�lW��S
����i�u��w�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�Ơ�lV��[��*ۊ�1�'�&�d�6�.��������@H�d��Uʹ�
�
�a�
������
�ד�@��Y1�����u�'�6�&��0�(�������P�������6�0�
��$�o�(���&���R��^	������
�!�d�1�0�E���Y����V��=N��U���u�3�}�4��2��������F�V�����&�$��
�#�l����K���G��d��U���u�u�u�9���Cځ�&¹��W��D_��Hʡ�%�l�
�0��m�N��T����\��XN�N���u�u�u�0�$�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����ԓ�@��G�����u�u�u�u�w�}�Wϲ�&ù��9��1�����&�u�h�4��2�����ғ�T�_�����:�e�n�u�w�}�Wϻ�
��ƹF�N��U���!�e�a�`�2�l��������[�o6�����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�#�m�C����ד�VV��D��ʥ�:�0�&�u�z�}�Wϲ�&ù��9��1��E���&�2�
�'�4�g��������C9��N��*���
�&�$���)�G���������D�����
��&�g��.�(��s���Q��Yd��U���u�<�u�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o�(���&���	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��G���8�g�|�|�w�5��ԜY���F�N��*ڊ�a�
�
�
�2�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�[��*��
�
�
�0�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�#�m�C����ד�VW��D��ʥ�:�0�&�u�z�}�Wϲ�&ù��9��1��D���&�2�
�'�4�g��������C9��N��*���
�&�$���)�E���������D�����
��&�g��.�(��s���Q��Yd��U���u�<�u�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o�(���&���	��F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��D���8�g�|�|�w�5��ԜY���F�N��*ڊ�a�
�
�
�2�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�[��*��
�
�
�0�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߊu�u�!�e�c�h���������h�����0�!�'� �$�:����5����2��x��G���3�
�b�m�'�t�\ϫ�
����WN��h��ۊ�;��;�0�6�9�4�������U�� ^�����n�_�u�u�z�1�(߁�Mƹ��9��N�����u�'�6�&�y�p�}���Y����lR��h��*���
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	���&����V�N�����;�u�u�u�w�4�W���Q����\��h�����u�u�%�6�~�<����	����@��X	��*���u�%�&�2�4�8�(���
����U��^��\���=�;�_�u�w�}�W���Y����lR��h��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W����֓�S��h_�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9F���*���
� �d�g��o�K�������T��A�����;�<�;�1�6�����&����lV�N�����0�}�
�0�"�)�B���&����l��UךU���4�
�
�
�"�l�@؁�K���@��[�����6�:�}�;�>�3�ǿ�&����G9��Z��\��� �&�2�0�������Г�F9�� ]��D���_�u�u�4���(���H����CU�
NךU���u�u�4�
�����NĹ����YN�����
�
� �d�d��D��Y���O��[�����u�u�u�
�2�(��������U��UךU���4�
�
� �f�o�(��E��ƹF�N�����
�
� �d�e��Eϩ�����@��h��*��g�e�u�u�f�t����Y���F������!�`�3�
�e�e���Y����V��[_�����c�f�%�u�j�W�W���Y�Ƣ�D5��1��*��m�%�u�=�9�u��������lT��1��]���h�r�r�u�;�8�}���Y���F*��C1�����!� �!�'��k�(ہ�����9��d��Uʻ�"�0�d�3��h�A���Y���F�N�� ���!��&�
�#�(����&����9��h\�M���u�=�;�}�2����&����W��G\��\��r�r�u�9�2�W�W���Y�ƹ�l��t��*��� �!�'�
�`��(���K����CW��N�����0�g�3�
�b�m����D���F�N��*����&�
�!�"�)����Oʹ��U��Y�����=�;�}�0��0�D�������N��S��D���0�&�u�u�w�}�Wϫ�&����R��d�����0�d�f�a�1��C���	��ƹF��R��ي� �g�m�
�d�a�W���Y�����d�����`�g�%�u�?�3�_�������U��X�����|�h�r�r�w�1��ԜY���F��@=��D���
�`�c�%�l�}�Wϰ�����l ��X�*��i�u�u�u�w�}��������V9��E�� ���d�c�`�3��i�O���Y����N��[1�����3�
�`�c�'�u�^��^���V
��d��U���u� �
�!��.�(�������V9��1�����a�m�%�n�w�}�����ӓ�F9��W��F��u�u�u�u�w�(�(���:����`��T����f�a�3�
�c�e�������@��C��B���
�`�c�%��t�J���^�Ʃ�@�N��U��� �
�!��$���������P��1��*��g�%�n�u�w�3� ���O����P��h�I���u�u�u�u�"�����
����A��B��D���`�3�
�a�o�-�W����ο�_9��G[�����`�e�%�}�~�`�P���Y����l�N��Uʠ�
�!��&��)�������� 9��Q��A���%�n�u�u�9�*��������S��N�U���u�u�u� ��)�4���&����P��R1�C���3�
�a�m�'�}����Q����G��h��*��e�e�u�u�f�t����Y���F������4�0��'�4�(���@�ғ�F9�� \��G�ߊu�u�0��;����J����Z�=N��U���u�0��9��(�E��&����[�������
� �g�c��o�G���Y�����RNךU���u�u�0��;����HĹ��l�N�����l�3�
�c�a�-�W��s���F�B"�����&�
�!� �#�/�(��&ǹ��lT��1��U���;�}�0�
�:�n����K����O�I�\ʰ�&�u�u�u�w�}��������V9��E�� ���d�c�`�3��i�O���B�����d�����`�g�%�u�j�W�W���Y�ƹ�l��t��*��� �!�'�
�a��(���K����CT��_��]���
�8�`�
�"�o�Cف�K���F�G�����_�u�u�u�w���������G��C��*��
�
� �g�a��F�ԜY�Ƣ�D��Y��*ۊ� �g�f�
�d�a�W����ԓ�9��h_�D���}�d�1�"�#�}�F��Y����V��P �����
�`�`�%�w�`��������U��W�����d�1�"�!�w�l�L���Yӈ��l��h��D���
�l�`�%�w�`�_���&����W��R�����3�
�l�a�'�}�Ϫ�	����]	��Q��L���%�|�_�u�w�2�(���&����U��^�����h�}�0�
�:�d�(�������l ��Z�*��:�u�8�
�n�3����&����l��d��Uʻ�!�=�g�3��n�(��E���F��R �����d�
� �`�f�-�W���	����@��AV��3���9�0�w�w�]�}�W�������U��W��G��u�e�u�=�9�u����N����Q��GZ��U���6�;�!�9�o��^ϻ�
���]ǻN�����&�
� �c�`�-�W��[����[����*���3�
�l�
�c�`��������_��q(�����u�d�n�u�w�3����&����
V��N�U��u�=�;�}�:��(���M�Г�F�V�����
�#�
��w�1����[���F��C��G���
�a�
�g�k�}�F������G��X�� ���d�%�u�u�'�>��������O��[��W���_�u�u�:�%�.�(���O�ӓ�F�L�U���;�}�8�
�o�;�(��&�����T�����g�
�|�0�$�}�G��Y����\��D[�� ��f�%�u�h�u�� ���Yے��lU��Q��Eߊ�d�h�4�
�8�.�(���J���V
��L�N���u�;�!�=��(�C���	���D�������8�
�
� �c�k����Y����\��h��F��u�9�0�w�u�W�W�������WW��B1�Bފ�g�i�u�&�;�)��������V��N��U���
�b�3�
�c�i����s���\��X ��*���g�l�
�g�k�}��������F9��^��Gʺ�u�'�6�;�f�;�(��M����l�N��*���1�d�<�
�"�o�Gہ�K�����hV�����e�m�%�u�9�}��������
T��G�U���:�
�:�1�f�4����O�ߓ�F�F����
� �d�d��o��������U��^�����_�u�u�'�4�3�N܁�H����W��h�I���!�%�m�
�"�o�Nׁ�KӇ����1��*��f�%�|�_�w�}��������Z9��h_�@���u�h�}�8��n����O�Փ�F��SN��ۊ� �d�c�
�e�f�W�������]��B1�Cڊ�g�i�u�&�;�)��������P��N��U���
�8�`�
�"�o�Eׁ�K��ƓF�C��*ڊ�0�
�9�=��-��������TF��D��U���6�&�{�x�]�}�W���&����R
��V1��*���
�;�&�2�6�.���������T��]���
�0�
�9�?������Ƽ�9��Q1�����4�
�9�
�%�:�}���Y����]l�N��Uʼ�u�}�%�6�9�)���������h��*���=�
�%�#�3�t����Y���F�N��U���
�0�
�9�?���������@��S��*ڊ�0�
�9�=��-����s���F�R��U���u�u�u�u�w�-�G�������[��G1�����
�<�u�h�'�m��������l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������_��h�����4�&�2�u�%�>���T���F��1�����%�4�<�
�>���������PF��G�����%�e�'�3�6�-����&ù��U9��G�����y�%�e�'�1�<��������WOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�e�'�3�6�-����&����F��R ��U���u�u�u�u�'�m��������l��D��I���
�
�0�
�;�5�L���Y�����RNךU���u�u�u�u����������Z��^	��Hʥ�e�'�3�4�'�<����B���F���U���u�u�u�0�3�-����
��ƹF��h_��&���:�u�h� ��.�4���&����P��R1�C���&�
�0�
�g�k�}���Y���C9��h=�����4�
�9�u�$�4�Ϯ�����F�=N��U���`��6�:��-��������]9��X��U���6�&�}�%�4�q��������V��c1��Gي�&�
�g�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���f�3�8�g�~�t����Y���F�N��U���`��6�:��-����E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���`��6�:��-����E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�H����l��h�����<�
�<�u�$�4�Ϯ�����F�=N��U���
�0�
�4��-��������T9��D��*���6�o�%�:�2�.��������R��G1�����
�
�0�
�6���������TOǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��%�d�'�3�:�%�������G��d��U���u�u�u�%�f�/��������E
��^ �����h�%�d�'�1�0����&����9F�N��U���0�_�u�u�w�}�W���&¹��U9��O1��*���
�;�&�2�k�}�(ށ�����K9��h��*���2�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����^��^ �����&�<�;�%�8�8����T�����h��*���
�;�&�2�6�.���������T��]���
�0�
�4�{�-�F�������l��PB��*ۊ�0�
�4�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h_�����4�
�%�#�3�t����Y���F�N��U���
�0�
�4��3����E�Ƽ�9��Q1���ߊu�u�u�u�;�8�}���Y���F�G1�����8�-�<�
�>�}�JϮ�H����l��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�x�w��(�������C9��S1��*���u�&�<�;�'�2����Y��ƹF��h\�����1�4�
�9��3��������]9��X��U���6�&�}�
��8��������WJ��h\�����1�4�
�9��/��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h\�����1�4�
�9�~�}����s���F�N������'�:�
�'�+����&����[��h\�����1�4�
�9�l�}�W���YӃ��VFǻN��U���u�u�
�
�2�4����&����Z��^	��Hʥ�g��'�:��-����	����9F�N��U���u�3�u�u�w�8�Ϯ�����lǑN��X���
�
�0�<�3�4�(���Y����T��E�����x�_�u�u����������@��V�����'�6�o�%�8�8�Ǯ�K����Z	����*���<�1�%�0�{�-�E�������R��[
��U���7�2�;�u�w�}�WϷ�Y�έ�l��D�����
�u�u�
��8��������WO�C��U���u�u�u�u�w�-�E�������Z��^	��Hʥ�g��'�:�l�}�W���YӃ��VFǻN��U���u�u�
�
�2�4����&����[��h\�����1�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�}�WϮ�M����Z��P1��E��u�!�
�:�>�����۔��Z��B �����}�!�e�a�b�8�G�������T9��^��F���n�_�u�u�z�-�C�������T9��1��*���u�&�<�;�'�2����Y��ƹF��hZ��*���<�2�0�e�6�����
����l��TN����0�&�4�
�2�}��������B9��h��F���8�g�|�u�w�?����Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�g�~�}����s���F�N������!�8�;���(������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�
�
�
�>�4����I����E
��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԜY�Ƽ�9��C�����
�u�h�6���2���+����lT��h��*���
�e�`�_�w�}�Z���&ǹ��G��Y	��*ۊ�%�#�1�4�$�:�W�������K��N������!�8�;���(�������@��Y1�����u�'�6�&��-�������T9��R��!���g�
�&�
�e�W�W�������F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�f�3�:�o�^�������9F�N��U���u�
�
�
�>�4����H����E
��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�%�c���������9��h��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C��*ߊ�0�
�0�4�6�����������^	�����0�&�u�x�w�}��������V��V�����;�&�2�4�$�:�(�������A	��D��*ߊ�0�
�0�4�6����	�ӓ�V ��R�����9�
�'�2�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l��h�����
�9�|�u�?�3�}���Y���F�G1�����7�!�
�%�!�9���������h��*���4�4�
�9�l�}�W���YӃ��VFǻN��U���u�u�
�
�2���������W9��h��U��%�`�'�3�5�)�(�������A��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�
�
�2���������TF��D��U���6�&�{�x�]�}�W���&����Q��h�����4�&�2�
�%�>�MϮ�������h��*���4�u�
�
�2�����	������h��*���4�4�
�9�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�Ƽ�9��Q1�����%�#�1�|�#�8�W���Y���F���*���
�0�4�<��4�W��	�ӓ�V ��R�����u�u�u�9�2�W�W���Y���F��1�����!�
�;�&�0�a�W���&����Q��h���ߊu�u�u�u�9�}����Y����]��E����_�u�u�
����������Z�D�����6�#�6�:��8��������]��[��*��
�
�
�e�{�o�^�ԶY���F��1�����;�
�
�
�'�+�Ͽ�
����C��R��U���u�u�%�c��)����&����R��[
�����;�%�:�u�w�/����Q����VJ��G1�����0�
��&�e�����K���F��P��U���u�u�<�u��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�D�������O��_�����u�u�u�u�w��(�������l��h�����i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϮ�O����Z��P1��E���
�9�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dךU���
�
�
�<�>�:���E�Ơ�lV��[��*ۊ�e�_�u�u�z�}�(ف�&����]��h_�����1�4�&�2�w�/����W���F�G1��7���8�;�
�
��-��������]9��X��U���6�&�}�%�4�q��������V��c1��Gي�&�
�g�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���f�3�8�g�~�t����Y���F�N��U���
�
�<�<�0�8�F���&����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�%�c��#�0����&¹��l��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��ԶY����l^��h:�����0�e�i�u�#�����&����\��R�� �&�2�0�}�#�m�C����֓�O�G����u�x�u�
����������l��A�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��c�����
�
�%�#�3�<����&����\��E�����%�6�y�4��4�(�������@��h��*��_�u�u�0�>�W�W���Y�ƥ�N�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C\�����g�|�|�!�2�}�W���Y���F��hV��*���<�2�0�e�6�����DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�������8�;���(������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�}�WϮ�A����Z��P1��D��u�!�e�a�b�8�F���B���F���*���<�<�2�0�f�<�(���Y����T��E�����x�_�u�u���(�������lW��G1�����&�2�
�'�4�g��������C9��N��*���
�&�$���)�D�������9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����T�N�����u�u�u�u�w�}����:����Z��R1�����9�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����p9��Z��*���
�%�#�1�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R�����u�%�l�
�f�;�(��I����[�e��ۊ�9�
�0�:�����Nƹ��	��E��*���g�`�
�g�l�}�WϮ�@ƹ��U��W�����h�}�4�2�f�<��������l ��X�*��:�u�0�d�1��B���	����F�G1�*���:�2�;�<��(�E��&���F��Z�����g�c�%�u�%�9��������\��h��G��
�f�n�u�w�-�N؁�����R��_�����3�
�f�l�'�}�J���&�ѓ�V��P��ۊ�0�
�e�e�/�/��������_��G�U���%�l�
�0�8�:��������T��N�U¡�%�
� �g�f��Eϱ�Y����G��M�����2�f�e�|�]�}�W���N����\��Y1�����3�
�f�l�'�}�J���&�ѓ�V��P�����
�f�g�%�w�2�W�������l
��h_����u�
�m�<��(�E��&���F��Z��F���
�d�d�%�w�3�W����ד�_
��R��*؊� �g�`�
�e�f�W���	����Z9��h_�L���u�h�}�8��h����O�ѓ�F��SN�����
�9�
�0�8����N����]ǻN��*��� �!�f�3��l�D���Y���^��a1�����e�f�%�u�9�}����Kù��lW�� 1��\�ߊu�u�
�0�"�)�B���&����l��S�����:�<�
�0�#�/�����ι�@��R
�����`�3�
�g�f�-�^��P��ƹF��h<�� ���c�3�
�e�d�-�W��
����\��h�����'�&�/�}�9�4��������9��h_�@���|�`�|�n�w�}����
����@9��h_�D���u�h�}�4�����K˹������*���3�
�f�`�'�t�}���Y����_T��h��D���
�g�c�%�w�`�}���Y���R��X ��*���g�����}����Q����T9��P1�L���|�h�r�r�w�1��ԜY���F��h�����#�g�e�_�w�}�(���K�֓�l��B1�Fߊ�f�i�u�u�w�}�WϿ�&����G9��\��3�����"�0�w�4����H����lT��F�U���d�|�0�&�w�}�W���YӇ��P	��C1��F؊�n�u�u�%��1�(�������W��N�U���u�u�u�!�'�k�(���H����CT��_��]���
�8�a�
�"�l�@ځ�K���F�G�����_�u�u�u�w�8�(���Jʹ��lW��1��N���u�%��9��o�G���@����K9��h\�E���u�h�_�u�w�}�W����ԓ�9��P1�G���=�;�}�'�2�:�(���J�ӓ�\��B1�Lފ�g�e�u�u�f�t����Y���F������!�9�f�
���1���s���C9��[\��G���<�8�-�3��n�F���Y���F�N�����9�
�
�0��d�@ϩ�����A��P��*���:�
� �g�d��E��Y���O��[�����u�u�u�%�4�3����J����u ��q(�U���%��9�
��(�F��&���FǻN��U���8�
�d�3��o�E���Y����N��G1�*���d�c�
�g�g�}�W��PӃ��VFǻN��U���
�4�g�e�>�4�(���H����CU��N�����9�
�
� �f�m�(��E�ƿ�W9��P�����:�}�;�<�9�9��������U��^�����~� �&�2�2�u����J����R��h�\�ߊu�u�
�4�e�i����M�ӓ� F�d��U���u�!�%�g��(�F��&����[����*���g�
� �d�o��E��Y���O��[�����u�u�u�0��0�Fց�����9��d��Uʥ��9�
�
�"�l�C؁�J���9F�N��U���
�d�
� �f�n�(��������h[�����m�e�%�}�~�`�P���Y����l�N��Uʥ��9�
�
�����Jƹ��l�N��#���
�
� �d�n��E��Y����_	��T1�����}�;�<�;�3�-�!���&˹��lW�� 1��\��� �&�2�0��0�(�������_��G����u�
�%�
�"�l�A܁�K���@��[�����6�:�}�;�>�3�Ǫ�	����l ��_�*��u�u�;�<�9�9��������_��G����u�
�%�3��m�@���Y����G��X	��*���!�'� �&�0�8�_���&�ד�F9��]��D���u�;�<�;�3�<�(���
����9��UךU���u�u�:�d�f�>��������9��R�����9�2�6�#�4�2�_�������Z��SF��ۊ�
� �g�d��o�[��P��ƹF��X��D���
�e�f�%�w�`��������l��C�� ���2�0�}�g�e�/���O�����^	��´�
�:�&�
�!�o�E���B���F���D���&�
� �d�d��F��Y����_	��T1�����}�0�<�0�$�:�����ד�F9��Y��G���g�|�_�u�w�-�ށ�����9��R�����9�2�6�#�4�2�_������� ��E��G��|�~� �&�0�8�_�������l
��1�\��u�u�u�u�'�.�(ށ�����F9��Y��D��u�!�
�:�>�����۔��Z��D�����:�g�d�3��m�E���P����]ǑN�����
�
� �g�e��E��Y����_	��T1�����}�;�<�;�3��(݁�����R�N�����0�}�%�6�9�)���&���l�N��Uʥ�&�
�4�!�1��B���	�����h�����0�!�'�'�$�'�_�������\��Q��@���%�|�f�|�l�W�W����ԓ�F9��X��G��u�!�
�:�>�����ۓ��Z��SF��*���
�l�f�u�w�3����ۇ��P	��C1��D؊�d�|�_�u�w�?�F���&����l��S��U���u�u�<�;�0�l����K����D��F����
� �d�`��o�G���Y�����RNךU���u�u�8�
�f�����@����F�F�����;�d�3�
�d�k����D�ξ�Z9��Q��F���%�u�;�u�5�;�(��@����l�N��*���<�;�f�3��e�D���Y���A9��^_�� ��b�
�g�4�3�,�(ށ�����9��UךU���7�3�
�f�n�-�W��s���F�^�����2�g�l�u�?�3�_���&�ғ�F9��Y��G��u�u�d�|�2�.�W���Y�����hY�����f�d�%�n�w�}��������S��N�U¼�8�f�3�
�f�l�����Ƹ�C9��h��D��
�g�n�u�w�/�!�������_��N�U���
�:�<�
�2�)�ǭ�����Z�������1�4�
�:�$�����J����u ��q(��3���:�<�!�2�%�(�������F�C��M؊� �g�d�
�f�n�Z�������V�G����u�
�
� �f�n�(��E�ƿ�W9��P�����:�}�=�3��4��������V��G1�����9�`�
����1���?���G	��Y�����;�<�;�1�p�z�QϪ�	����U��\�����d�d�1�"�#�}�^���P���F��Q��F���%�u�h�}�4�-�(���&��������*���3�
�f�b�'�t�}���Y����ZW��B1�BҊ�g�i�u�!�'�l�D���&����l��X��*ۊ�0�
�l�g�l�}�WϬ�����F9��^��G��u�!�%�d�e�;�(��O����\��h��D��
�g�n�u�w�/�ށ�����9��R��]���
�e�
� �f�h�(������C9��Y�����d�n�u�u�%�+�(���H����CT�
N�����e�
� �d�n��DϦ�Ӈ��P	��C1��D��n�u�u�'�!����L����Z���*��
� �g�a��n��������]��[��D��u�u�'�#��(�E��&���F��Z��GҊ� �g�m�
�d�%�Ͽ�&����G9��1�N���u�'�#�3��j�(��E����\	��O)��:����0�!�'������&����T9��\�����%�6�;�!�;�l�F��Y����V
��Z�*���m�l�%�u�j�W�W���Y�ƿ�_9��G[�� ��`�%�u�=�9�u����M����_��G\��\��r�r�u�9�2�W�W���Y�ƹ�l��t��*��� �!�'�
��(�@���	��ƹF��R����
� �l�b�'�}�J�ԜY���F��h�����#�
�u�=�9�u�����Փ�F9��1��]���h�r�r�u�;�8�}���Y���R��X ��*���
�n�u�u�$�1����K����R��h�I���u�u�u�u�#�-�A؁�����9�������8�
�`�'�0�o�E���P���A�R��U���u�u�u�4��2�����ԓ�l�N�����%�f�1�8�%�<�(���N�ߓ�F�F�����%�
�0�:�0�3����Mʹ��	��C��G���
�m�
�g�l�}�Wϭ�����U��B1�Fي�g�i�u�!�'�l�(���&�����������!�9�d�d�l�}�Wϭ�����R��B1�FҊ�g�i�u�!�'�l�(���H����CT��Y
�����8�d�
� �f�n�(��B�����h��D���1�8�'�4��(�F��&���F��Z��C���2�g�b�u�%�)���&����Q��G\����u�0�
�8�f����Mǹ��Z���*���d�
� �d�d��EϿ�Ӓ��l_��Q��F���%�|�_�u�w�8�(���HŹ��lW��1��U��_�u�u�u�w�����J����R��h����u�&�9�!�'�h����M�ғ�N��S��D���0�&�u�u�w�}�Wϭ�����T��B1�G܊�f�_�u�u�2����&����S��G\��H���8�
�l�3��n�O���Y����R��X ��*���
�|�_�u�w�8�(���H˹��lW��1��U��}�0�
�8�f����J˹������*���d�
� �d�b��E��Y����V
��Z�M���8�'�4�
�"�o�Fف�K�����hV�����a�a�%�u�%�)���&����^��G\����u�0�
�8�f����Nù��Z�=N��U���u�
�4�g�d�;�(��O����D��F�����%�m�3�
�c�i����P���A�R��U���u�u�u�&�;�)��������V��UךU���0�
�8�d�1��D߁�K�����G1��*��
�g�-�'�6�����&����O��N�����!�%�e�
�2�2�������� R��N�U¦�9�!�%�l��8��������S��h����8�
�e�3��i�C���P���F��[1�����3�
�a�f�'�}�J�������C_��S�����
� �d�b��o��������]��[��D��u�u�&�9�#�-�F���&����l��S�����m�3�
�g�a�-�W���Y����G��1��*��f�%�|�_�w�}��������U�� ^�����h�}�8�
�g����Lʹ��	��C��Aي�:�
� �d�g��E��Y����V
��Z�*���d�d�
�g�k�}����MĹ��lW��1��U���u�0�
�8�e����Iʹ��]ǻN�����8�g�
� �f�o�(��E��ƹF�N�����d�4�9�:�2��(���H����CT��_��]���
�8�g�
�"�l�Fځ�K���F�G�����_�u�u�u�w�8�F���&����l��=N��U���
�8�g�
�"�l�D؁�J���9F�N��U���2�d�4�9�-�/����&����l��@��U¦�9�!�%�f�1��@���	����[�I�����u�u�u�u�w�-�Nځ�&����_��G\�U���&�9�!�%�a�;�(��N����[�C��F݊� �d�`�
�e�%�Ͽ�&����G9��1�N���u�&�9�!�'�j����J�ԓ�F�F��؊�0�
�e�f�6�9��������lT��G�U���&�9�!�%�o�;�(��O����[�C��F݊�0�
�e�f�6�9��������lT��G�U���&�9�!�%�n�;�(��J����[�N��U���4�
�:�&��+�E��������hX�����f�m�%�}�~�`�P���Y����l�N��Uʥ��9�
�
�2��N��s���@��C��*���b�c�%�u�j�u��������l��V �����!�%�
� �`�m����s���@��C��E���
�f�e�%�w�`�_���&�ד�V��^����4�
�:�&��+�(���s���@��C��D���
�f�`�%�w�`�_�������U��Z�����;�u�0�
�:�n�(���K����CT�=N��U���
�8�f�
�"�l�F܁�J���9F�N��U���
�d�
�0��d�Fϩ�����^��1����b�}�|�h�p�z�W������F�N��*���&�
�#�g�g�W�W�������CU��Q��L���%�u�h�}�:��A�������F��EN��*���&�
�#�
�~�W�W�������CU��Q��L���%�u�h�}�:��D���&����l��V �����!�%�f�3��d�N���P���F��[1�����3�
�l�e�'�}�J�������CU��Q��L���%�u�;�u�:��E݁�����9��UךU���0�
�8�f��(�F��&���FǻN��U���
�4�g�l�1��O���	�ƻ�V�D�����`�3�
�l�g�-�_���D����F��D��U���u�u�&�9�#�-�E���&����l��=N��U���
�8�f�
�"�l�Cہ�K�����h_�*���d�c�
�f�/�/��������_��G�U���&�9�!�%�o�;�(��I����[�D�����a�3�
�l�c�-�W���Y����G�� 1��*��a�%�|�_�w�}��������U��[�����h�_�u�u�w�}�(���K�ߓ�F9��]��Gʢ�0�u�&�9�#�-�O���&����l��G��U��|�0�&�u�w�}�W���
����^��h��D��
�f�_�u�w�8�(���J����_��G\��H���8�
�
� �a�m�����ƿ�_9��G1��*��
�g�n�u�w�.����	�֓�F9��W��G��u�&�9�!�'�h�(�������l ��W�*��-�'�4�
�8�.�(���&����F�D�����d�3�
�l�b�-�W��Q����9��h_�C���u�;�u�0��0�C߁�����
9��UךU���0�
�8�a��(�E��&���F��Z��G܊� �g�a�
�d�2�W���&�֓�\��B1�M܊�g�n�u�u�$�1����J����W��h�I���!�%�m�
�"�o�Aց�KӇ����h��A؊� �g�l�
�e�f�W���
����^��h��G��
�f�i�u�w�}�W���+����9��[1�����
� �g�b��o� ���Yە��l��]�� ��l�
�g�e�w�}�F�������9F�N��U���f�3�
�e�d�-�L���Yӕ��l��[�� ��g�
�f�i�w�}�W���YӴ��T��V�����&�g�3�
�f�j�������@��C��F���
�d�m�%��t�J���^�Ʃ�@�N��U���%�l�
�d�1��F���	��ƹF��R����
� �g�`��o�K�������9��h\�L���u�:�u�%�4�3����H���9F���*���a�
� �g�a��E��Yے��9��h\�G���u�;�u�&�2��(���&����]ǻN�����8�a�
� �e�j�(��E����^��1��*��l�%�u�;�w�.����&����_��UךU���0�
�8�a��(�E��&���FǻN��U���%�6�;�!�;�n�(������G��Y�� ��d�
�g�e�w�}�F�������9F�N��U���4�g�d�
�2��G��s���@��C��*���m�g�%�u�j�W�W���Y�ƪ�l'��O!��*���:� �0��;�8�N؁�����T��_��]���
�8�b�3��k�(��I���W����ߊu�u�u�u�2���������9��d��Uʦ�9�!�%�e�1��C���	���N��G1�*���
�l�m�-�%�<�(���
����9��d��Uʦ�9�!�%�d�1��C���	���N��Z��ۊ� �g�e�
�e�<�ϭ�����V��B1�GҊ�g�n�u�u�$�1����K����S��h�I���!�%�m�
�"�o�Oہ�KӞ����T�����d�d�n�u�w�.����	�Փ�F9��^��G��u�!�%�m��(�E��&����]��R�����
� �g�e��o�L���Yӕ��l��Z�� ��g�
�g�i�w�.����	����W��E	��*���g�d�
�g�/�/��������_��G�U���&�9�!�%�b�;�(��A����[�C��Lڊ� �g�l�
�e�<�ϭ�����R��B1�G؊�g�n�u�u�$�1����O����S��h�I���&�9�!�%�g���������F9��Z��Gʭ�'�4�
�:�$��ށ�P���F��[1�����3�
�`�c�'�}�J�������l ��Z�*��4�1�&�9�#�-�A���&����l��d��Uʦ�9�!�%�
�"�e�B���Y���F�N�����:�&�
�#��}����Q����G��h��B���%�}�|�h�p�z�W������F�N��*���&�
�#�
�l�}�Wϭ�����9��Z����� �b�l�%�w�`�_���	����Q��G\��ʧ�#�3�
�b��o�L���Yӕ��l��1��*��
�g�i�u�5�2�(��� ����t��C��:���$�4�
�
�2��O������P��Y�����`�
�g�n�w�}��������U��X��G��u�!�%�g�1��Oہ�KӇ����h��C���
�c�
�g�l�}�Wϭ�����9��hV�*��i�u�u�u�w�}��������V9��E�� ���f�
�
�0��j�Oϩ�����P��Q��Bي�g�e�u�u�f�t����Y���F������4�0��'�4�(���&����^��UךU���0�
�8�l��8��������R��h�I���!�%�d�
�2��N���Ƹ�C9��h��D��
�g�n�u�w�.����	ʹ��l^��h�I���u�u�u�u�1�����
����A��B��Fۊ�
�0�
�b�o�*����
����^��Q��F܊�g�e�u�u�f�t����Y���F���*���m�3�
�g��n�}���Y����G��Q��Mߊ�g�i�u�&�;�)��������T��Q��Bӊ�g�-�'�4��2����¹��l�N��ۊ� �d�m�
�e�a�Wǲ�&����^��G_�����0�d�3�
�b�j����s���G��h��D��
�g�i�u�9�*��������lW��1��U���u�0�
�8�e����OĹ��]ǻN�����3�
�f�m�'�}�J���
����A��V�U���&�9�!�%�a�/���H����F�C��*���g�e�
�g�k�}����
����^��Q��L���%�u�;�u�:��C���&����l��d��Uʡ�%�
� �g�`��E��Yۊ��9��h\�M���u�;�u�0�d�;�(��J����l�N��܊� �g�c�
�e�a�Wǰ�����Q��1��*��d�%�u�;�w�8�(���MŹ��lT��1��\�ߊu�u�8�b�1��E���	���N��Y��D���2�g�a�u�%�.����	�Г�F9��X��G��u�u�!�%��(�E��&���F��S1�����#�6�:�}�9�4��������)��h\�*���4�
�
� �e�n�(��Y�ƹ�@��R
��*؊�0�<�1�<��4�^��Y����^��\�� ��m�
�d�i�w�����K����U��h�D���d�1�"�!�w�t�}���Y����V��Q��A���%�u�h�%��1�(܁�����9��]����!�u�d�n�w�}����H�ӓ�F9��W��F��u�:�d�3��h�@���Q����\��XN�\�ߊu�u�8�
�g����@ʹ��Z�G��*���d�f�
�g�f�}��������l�N����m�3�
�e�b�-�W������e9��Q��E���%�}�f�x�f�9� ���Y����F�C��Dڊ� �c�b�%�w�`�_Ǽ�����v��C1�����'��
�$�6��(���&����@��E�� ��g�%�|�s�0�-����MĹ��]ǻN�����d�
� �d�a��F��Y����l0��h��D��
�d�`�u�w�}�������9F���*��
� �d�e��l�K�������9��h_�F���}�g�x�d�3�*����P���F��G1�G���
�m�c�%�w�`�1݁�&����^��G]��Dʱ�"�!�u�|�]�}�W���&����U��]�����h�!�%�c��(�F��&���F�N�����u�|�_�u�w�0�(��&����T��G]��Hʸ�;��c�3��m�D���Q����]��R�����;�1�!�%�a���������_��G�����!�u�:�<�#�:�ǫ�
����WN��G1�*���!�3�
�d�n�-�^���������^ ����� �&�2�0��0�(�������U��_�����k�u�u�;�w�2��������]��Y�����c�
�4�!�1��F���	���S�������w�_�u�u�:��Fځ�����9��R��3؊�
� �d�l��o�F�������W�=N��U���
�d�
� �f�h�(��E�Ƹ�C9��h��D��
�g�c�x�f�9� ���Y����F�C��D���3�
�d�l�'�}�J�ԜY���F��h�����#�
�c�"�2�}����Nù��lW��1��]���h�r�r�u�;�8�}���Y���C9��1��*��f�%�n�u�w�)���A����W��h�I���!�
�:�<��8��������VN��D�����8�
�d�
�"�l�Aց�J����O��N�����d�l�3�
�f�l����Dӕ��l
��^�����'�&�<�!�;�;�_���������T�����`�
�����1���?�ʸ�l��R	��]���<�;�1�r�p�{����H�ޓ�F9�� Y��D��x�u�:�;�8�m�^���B�����h_�����c�
�g�i�w�l�W����θ�C9��h��L���%�u�u�%�4�3����O������RN��W�ߊu�u�8�
�e����AĹ��Z���*��
� �d�m��o��������]��[�*ٓ�������L���YӒ��lW��h��D��
�f�i�u��<�E�������Q��F�U���;�:�f�|�]�}�W���&����U��Y�����h�%��9�����MĹ��W�_�����:�e�n�u�w�)���M����^��h�I���
�4�g�l�1��O���	������Y��F���_�u�u�8��o�(���K����CU�
N��ۊ�
� �g�d��o�F�������W��d��Uʡ�%�d�m�3��m�C���Y����\��1��*��g�%�}�d�3�*����H��ƹF��Z��G���
�g�
�a�k�}�$���&����l5��B�����g�!�
�;��(�B���	������Y��G���_�u�u�8��n����K�ӓ�F�L�U���;�}�<�;�3��(���&����F�D�����%�6�;�!�;�l�(���Y����D��d��Uʡ�%�d�
� �f�i�(��E�ƿ�W9��P�����:�}�;�<�9�9��������_��h^��Xʠ�&�2�0�}�e�/���H���9F���*���3�
�b�
�e�a�W��Y����N��G1�����3�
�a�
�c�`��������_��hZ�\ʰ�&�u�e�n�w�}����HŹ��lS��h�I����6�
�4�2���������9��h��*���`�b�%�}�d�p�FϺ�����O��N�����d�
� �d�a��E��Y���D��F�����0�}�g�a�1��E���	�����^	��´�
�:�&�
�!�o�D���Y����D��d��Uʡ�%�d�
� �b�j����D�΢�G��1��*��
�g�:�u�8�1�݁�����l��d��Uʡ�%�d�
�:��(�F��&���F��T��*���d�b�
�g�/�/��������_��G�U���!�%�d�3��e�(��E�ƪ�l��t��*��� �!�'�
�e�)�(���&����U��F�U���u�:�;�:�g�f�W�������9��h_�G���u�h�&�1�;�:��������A��M�����;�1��
��<����&����l��[�\�ߊu�u�8�
�f�;�(��O����[��C
�����
�0�!�'�$�4��������Z��SF�����3�
�g�m�'�t��������AN��D�����e�u�u�8��m����K�ԓ�N��_�����:�e�|�|�l�}�WϪ�	����U��^�����h�&�1�9�0�>�����ο�Z ��[��]���<�;�1�!�'�k�(���H����CW�C�����0�}�;�<�9�9�P���_Ӡ��9��D�� ��`�
�d�f�z�}�������O�=N��U���
�a�3�
�d�j����D������YN�����1��
�0��d�D���Y����V��G1�����9�d�
�c�~�8����I��ƹF�N�����`�6�&�
�"�l�E؁�H���@��[�����6�:�}�0�>�8�����θ�C9��h��D��
�g�y�g�~�W�W�������9��h_�G���u�h�&�1�;�:��������F��P ��]���'�2�g�d�~�v��������R��X ��*���g���|�]�}�W���&�ѓ�F9�� 1��U��3�
�!��$���������Q��X1�����
�b�
�d�d�}��������l�N����
� �`�b�'�}�Jϸ�&����R��d�����0�g�
�:�>�)����N����T��N����!�u�|�_�w�}����@����V��h�I���!�
�:�<��8��������]��q\�� ��f�%�|�~�"�.����Q����\��h��G����|�_�u�w�0�(݁�����l��S��D���=�;�}�8��m����LĹ��[��G1�����9�f�`�u�;�8�U���s���G��^�� ��e�
�g�i�w�l�W����ο�T����*���3�
�e�d�'�t�Iϭ�����R��X ��*���g�f�|�u�;�8�U���s���G��_�� ���`�%�u�h�1��5�������@	��C�����
�
�:�3��d�(��J�ƨ�D��\�N���u�!�%�f��(�F��&���F�N�����%��&�9�����O¹��[��G1�����9�`�
�|�2�.�W��B�����h]�����a�g�%�u�j�.��������V��EF�����}�;�<�;�3�,�(�������l ��]�*��y�g�|�_�w�}����M����V��G_��Hʳ�
��-� ��?��������F��h�����l�
�d�g�w�}�W������]ǻN�����`�3�
�g�f�-�W��Q����\��h��*���u�8�
�f�%�:�E��P���F��G1�*���d�g�
�g�k�}����H�Փ�F9��\��Fʭ�'�4�
�:�$��ށ�P���F��G1�*���d�`�
�g�k�}�F������@��R
�����3�
�`�b�'�t�Kϭ�����R��X ��*���g�f�|�u�;�8�U���s���G��V�� ��d�%�u�h��2����&����S��N��U���9�&�
� �a�d����s���G��W�� ��b�
�d�i�w�)�(�������P������� �&�2�0��2�F���
����lW��1��\���|�n�u�u�#�-�D���&����CR�
N��*����&�
�!�"�)����K����Z��Q��Cي�d�f�u�:�9�2�E���s���G��^�� ��b�
�g�i�w�)�(�������P�������<�=�}�<�9�9����/����T��h�Y���<�!�2�'�"�.����Q���F��G1�*���d�b�
�d�d�p�W������O�UךU���8�
�d�3��n�(��E����\��D[�� ��f�%�u�'�9�)��������9��UךU���8�
�g�3��i�(��E����^��1��*��
�g�4�1�#�-�Cށ�����l��d��Uʡ�%�a�
� �f�l�(��E���F��R �����0�}�:�g�1��B���	�����Y�����:�&�
�#�e�n�^������D��N�����a�
�:�
�"�l�G܁�K�����hZ�����c�f�%�u�8�}��������EW��UךU���8�
�a�3��k�B���Y����G��X	��*���!�'�'�&�-�u��������\��T��*���d�a�
�d�{�i�^�ԜY�Ƹ�C9��h��D��
�g�i�u�f�}����Q����VT��h_�� ��g�
�g�h�6�����&����lV�R��U��n�u�u�!�'�i�(���M�Փ�C��RN�U���6�;�!�9�b�n�}���Y����P��B1�F���u�h�3�
�#���������F��Y�� ���l�%�n�u�w�)���&����U��N�U������!��.����&����V9��h\�� ���a�%�n�u�w�)���&����^��G\��H���w�"�0�u�'�.�(���H����CT������!�9�d�
�a�}����[����F�C��AҊ� �g�l�
�e�a�Wǌ�����R
��X ��*؊�
�d�'�2�d�l�W���Y����\��h��*���_�u�u�8��d����I�ѓ�F���*���<�
�0�!�%�/����Q����T����*���
�
�
� �f�i�(��U���l�N�����3�
�l�
�e�a�W��Y����N��G1�*���c�b�%�u�w�-��������lP�R��U��n�u�u�!�'�h�(���H����CU�
N�����;�!�9�d�f�{����H�֓�F9��_��D��u�u�!�%�b����@¹��Z�_�����u�!�%�d�o�;�(��L����F��h�����#�f�e�u�;�8�U���s���G��\�� ��c�%�u�h��2����<����l!��V��*���� �9�&�%�:�E��Y�ƫ�C9��hZ�*��n�u�u�!�'�h�(���H����CT�
N��Wʢ�0�u�&�2�2�u�E�������
P��P�����1�4�
�:�$�����I����_��^�����u�8�
�a�1��N܁�K�����h��G���
�f�
�g�8�}�������� 9��UךU���8�
�`�3��j�C���Y����G��X	��*���!�'� �&�0�8�_�������l
��1�U���;�<�;�1���(���&����O��N�����`�
� �d�g��E��Y���D��F�����%��d�3��m�@���Y�ƭ�l��D�����a�f�u�9�2��U�ԜY�Ƹ�C9��h��L���%�u�h�}�2���������9�������!�%�
� �`�k����s���G��V�� ��e�
�g�i�w�l�W����ι�@��R
��G���3�
�b�l�'�t�Kϫ�
����WN��h�����#�g�f�|�w�1����[���F��G1�*���l�b�%�u�j�4����&���� U��F�U���u�:�;�:�g�f�W�������9��h\�M���u�h�}�8��l����K����\��Y
�����
� �g�d��n�L���YӒ��lP��Q��M���%�u�h�&�3�1��������AN��D��]���<�;�1�����������
P��G�A���_�u�u�8��l��������_��N�U¼�8�g�3�
�o�k�����ƭ�l��D��ۊ�|�_�u�u�:��E���&����l��S�����:�<�
�0�#�/��������[��^	��¸�;��c�'�0�o�B�������G��EF�����0�}�e�u�w�0�(�������T��F�X���:�;�:�e�~�t�L���YӒ��lP��Q��Cي�d�i�u�'�0�����J����S��N����!�u�|�_�w�}����M����^��h�I���!�
�:�<��8����
����l
��CF�����0�}�8�
�f�����@���G	��Y�����;�<�;�1�p�z�QϘ�&ƹ��@��B1�L܊�d�f�x�u�8�3���P���9F���*���3�
�m�`�'�}�J���[ӑ��]F��^	���
�
�0�
�n�i�W���������T�����d�
�c�|�2�.�W��B�����hX�����d�f�%�u�j�.��������V��EF�����0�}�g�g�1��G���	�����^	��´�
�:�&�
�!�o�1���P���F�N����
�4�!�3��l�N���Y����G��X	��*���!�'�'�&�-�u����ے��lP��Q��D���%�|�f�|�l�W�W�������l ��\�*��i�u�4�
��(�F��&���F�N�����u�|�_�u�w�0�(�������Q��N�U���
�:�<�
�2�)�ǫ�
����WN��h\�� ��l�
�g�u�w�3����ۇ��P	��C1��D؊��|�n�u�w�)���&����P��GZ��Hʓ�
�
� �d�c��D��Y����G	�UךU���8�
�
� �a�k����D������YN�����e�3�
�`��i�JϿ�&����G9��1�U���0�w�w�_�w�}����I����W��h�I���d�u�=�;��4��������9��h_�B���|�k�&�2�2�u��������EW��[��U���0�w�w�_�w�}����H����T��h�I���8�
�d�3��o�A���Q���W��X����n�u�u�!�'�j�(���H����CT�
N��Wʢ�0�u�%��$�1�(܁����� 9��S�����;�!�9�`��t����Y���9F���*���3�
�m�l�'�}�Jϭ�����Z��R��§�&�/�}�;�>�3�ǯ�&����T��h��D��
�g�y�g�~�W�W�������l ��W�*��i�u�!�%�f�i����A�ߓ� F��EN��*���&�
�#�
�~�W�W�������l ��^�*��i�u�d�u�?�3�_�������\��1��*��f�%�|�i�$�:����	����@��A_��F���u�9�0�w�u�W�W�������l ��]�*��i�u�4�
��(�F��&����\9��C�� �&�2�0�}�:��B���
����lW�� 1��\���:�;�:�!��3����Q����T����*���6�&�
� �f�o�(��P�ƻ�V�C�����0�}�;�<�9�9����Kƹ��@��B1�G݊�d�|�h�e�6�9��������AN��D�����8�
�`�6�$����KĹ��O�]�����u�x�n�u�w�)���&����S��G_��Hʦ�1�9�2�6�!�>����������^	��¥�&�
�
�4�#�;�(��A����S��UךU���8�
�m�3��m�D���Y����G��X	��*���!�'�&�<�#�/����
����WN��Y1��C���2�g�`�|�#������ι�@��R
��E���u�8�
�b�1��G���	����W��X����|�|�n�u�w�)���&����S��N�U���3�
�b�
�e�l�W������]ǻN�����e�3�
�e�o�-�W��[����[�������%�&�
�
�"�o�E݁�K���@��R
�����;�!�9�d��k�^ϻ�
���]ǻN�����e�;�!�3��l�A���Y���G��^�� ��l�
�g�-�%�<�(���
����9��d��Uʡ�%�m�
� �f�l�(��E�Ƹ�C9��h��D��
�g�c�x�f�9� ���Y����F�C��M؊� �g�d�
�f�a�W���&����P9��T��]���<�0� �&�0�8�_���K�ד�R��Q��E���%�|�`�|�l�}�WϪ�	����U��[�����h�w�w�"�2�}�%������� 9��h\�A���u�u�%�6�9�)���&����_��^�����u�8�
�a�1��G���	���l�N��Uʴ�
�:�&�
�!��Aϩ�����^��1��*��b�%�}�|�j�z�P������F�N�����
� �d�d��o�}���Y����S��B1�Cӊ�g�i�u�d�w�5�����ԓ�l ��^�*��h�4�
�:�$�����J����_��^�����u�8�
�c�1��E���	���N��Y	��*���
�;�&�g�>��E���&����l��O�����:�&�
�#��t�}���Y����Q��B1�Mފ�g�i�u�d�w�5����;����p��h=�� ���'�
�a�
�2��O��DӇ��P	��C1��F���u�9�0�w�u�W�W�������l ��Z�*��i�u�d�u�?�3�_�������@��C�����
�a�
�0��e�@������]��[��G���9�0�w�w�]�}�W���&�ߓ�F9��X��D��u�!�
�:�>�����۔��Z��B �����}�8�
�a�%�:�E��P����]ǻN�����
� �`�g�'�}�J�������l ��W�����'�;�!�=��(�C���	����F�C��Lڊ� �g�l�
�e�a�W��Y����N��h��6���
�!� �!�%��Cف�����Q������!�9�f�a�w�1����[���F��G1�*���g�l�
�g�k�}�F������F$��D1�����!� �!�'��i�(���&����[��G1�����9�f�c�u�;�8�U���s���G��]�� ��l�
�d�i�w�)�(�������P������� �&�2�0����������\��h��*��|�c�|�n�w�}����@ǹ��lW��1��U��&�1�9�2�4�+����Q����G9��Q�����;�1�4�
�8�.�(���M�Պ�u ��q(��3���y�:�<�!�0�/��������V�N����
� �d�a��l�D��Y����G	�G��\�ߊu�u�8�
�b�;�(��I����[�L�����}�;�<�;�3�?����H����BV�N�����0�}�
�
�2�4����&����F��D��E��u�u�!�%�n����Lƹ��Z���*���3�
�f�l�'�}����	����@��A[��F��������t�}���Y����
Q��B1�D݊�g�i�u�!�'�h�(���&����	��B �����"�d�'�2�d�n�^�ԜY�Ƹ�C9��h��D��
�f�i�u��<�E�������_��F�U���;�:�f�|�]�}�W���&����W��G\��H���:�
�0�
�:����Iʹ������*���3�
�a�e�'�t�}���Y����@9��hW�*��i�u�!�
�8�4�(�������V��RF�����0�}�-�
�:��(���@�ߓ�O�G����u��6�
�6�8�$�������lW��h�����
�c�e�%�w�`��������l��C�����/�}�;�<�9�9����
����V9��E�� ���d�c�'�2�e�h�^��P���F��h��6���
�!� �!�%��Cف�����l��S��U���u�u�&�9�#�-�F���&����CU��_��]���
�b�3�
�f��E��Y���O��[�����u�u�u�0��0�F߁�����l��=N��U���6�
�4�0��/��������F9��1��U��_�u�u�u�w�-��������lW��_��]���
�
� �c�a�-�_���D����F��D��U���u�u�4�
�8�.�(���&��ƹF��{1��*���0��'�6�"�8�F���M����R��h�I���!�
�:�<��8��������]��B"�����&�
�!� �#�/�(��&ƹ��lT��1��\��� �&�2�0����������9��T��#���
�f�d�%�~�f�W�������l%��R1����� �0�d�l�1��A���	���l�N��Uʻ�"�0�f�3��h�@���Y����N��h��؊� �g�l�
�e�m�W���H����_��=N��U���u�0��9��(�E��&����F�B"�����&�
�!� �#�/�(��&¹��lT��1��U�� �
�:�0�#�/�(��&����S��G\��Dʱ�"�!�u�|�]�}�W�������@��C�����
�b�
�
�"�o�Aׁ�H���@��[�����6�:�}�0�>�8��������F*��C1�����!� �!�'��j�(ށ�����9��B�\��u�u� �
�#���������F��Y�����c�e�%�u�j�W�W���Y�Ƣ�D5��1��*��g�%�u�=�9�u�����ԓ�F9��[��G��u�u�d�|�2�.�W���Y�����d��*���g�g�
�f�]�}�W�������@��C�����
�m�
�
�"�o�@ׁ�K���@��[�����6�:�}�;�>�3�ǫ�&����R��d�����0�d�l�a�1��C���	�����^	�� �
�f��!�e�i��������F9��W��F���_�u�u��4�����*����G��h_�*���g�b�
�f�k�}�W���Y����V��[_�����c�f�%�u�?�3�_�������l ��[�*��e�u�u�d�~�8����Y���F��R��ӊ� �g�`�
�d�W�W���5����V9��E��GҊ� �g�`�
�e�a�W���&����P9��T��]���<�;�1�!�'����MĹ��F�B �����}�� �g�"��D݁�����e9��h\�D���|�n�u�u�"�����&����R��h��*���'�0�g�3��j�B���Y���F�N�����e�d�a�
�g�*��������9��h\�E���}�|�h�r�p�}����s���F�G1��%���:�
�;�&�0�W�W���5����|��]�����9��3�
�d�l����D���F�N��#���
�g�e�<�:�%����J�ד� F��R �����!�%�d�3��n�B���Q���A��N�����u�u�u�u�$�1����@����U��h����u�� �g�"��Dہ�����e9��h\�L���u�h�_�u�w�}�W����ԓ�9��^\�*���
� �g�d��n� ���Yە��l��_�� ��f�
�g�e�w�}�F�������9F�N��U���
�8�a�
�"�o�Eށ�J���F��h��9����!�g�`�1��@���	�����h�����0�!�'�'�$�'�_���������O#��!ػ� �
�
� �e�l�(��U���l�N��*����g��!�$�;�(��N����[��{1�� ��� �
�d�
�"�o�F݁�K����W	��C��\�ߊu�u��-��$����H����lT��1��U��&�1�9�2�4�+����Q����T����*���<�1�<�
�>�t�Zϫ�
����WN��h��ۊ�;��;�0�6�9�4�������U�� ^�����n�u�u� �3�/����H����T��h�I���u�u�u�u�#�-�Oف�����9�������0�
�8�a��(�E��&���F�_��U���0�_�u�u�w�}��������U��X����u�u� �1�%�1� �������F9��W��G��u� �1�'�;�*�F�������F��EN��*���&�
�#�
�~�W�W�������_	��Q��F���%�u�h�_�w�}�W�������l ��\�*��"�0�u�&�;�)��������P��F�U���d�|�0�&�w�}�W���Yӕ��l��Y�� ��e�
�g�_�w�}��������]	��Q��F���%�u�h�}�9�8����&���� W��G]�����%�6�;�!�;�l�F������V��d