-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�e�����}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e��o��w�	�(���0����p2��F�U���;�:�e�n�w�}��������}F��s1��2���_�u�u�
����������}F��s1��2���_�u�u�
��<�W���7ӵ��l*��~-��0����}�d�1� �)�W���s���C9��Z�����9�u�u����;���:���F��1�����u�u�����0���/����aF�N�����u�|�_�u�w��(�������C9��SN�<����
���l�}�WϮ�M����Z��P1��E��������4���:����U��S�����|�_�u�u���(�������lV��G1����������4�ԜY�Ƽ�9��c�����
�u�u� �w�	�(���0����p2��F�U���;�:�e�n�w�}����,����Z��R1�����9�u�u� �w�	�(���0��ƹF��h[��U���������!���6���F��@ ��U���_�u�u�
����������}F��s1��2���_�u�u�
����������\��b:��!�����
����_������\F��d��Uʥ�c���8�9��(߁�	����\��b:��!�����n�u�w�-�A���-����T9��N�:���������4���Y����W	��C��\�ߊu�u�
�
��4�����ד�C9��SN�:��������W�W���&Ĺ��	F��=��*����
����u�FϺ�����O��N������4�
�9�w�}�9ύ�=����z%��N������!�8�;���W���,�Ɵ�w9��p'��#����u�f�u�8�3���B�����h9�����2�0�e�4��1�W���,�Ɵ�w9��p'�����u�
�
�
�>�4����H����f2��c*��:���
�����l��������l�N��M���!�8�;�
����������f2��c*��:���n�u�u�%�f���������f2��c*��:���
�����}�������9F���@���6�:�
�%�!�9�Mϑ�-ӵ��l*��~-��N��1�_�_�'�?�)����ӄ��R��QN��Eߔ���
�u�$�W�W�������F��t!��*���������W���-����l�N����� �0�����2���0����} ��X�����u�u�'�=�#�>�������F��r^��B���3�e�=�&�>��G���Mߝ��`9��g;��!���h�-�y����"���5����J��d1��%������e���>���-����g[�� �E���a�a�d����'���:����T��^�E����
�� ���?ұ�����{*��d7��6����g�{�b�g�m�?���*����r2�B��&������;�9�q�;��� ����~[��"��&�����g�y���.���?����J��d1��;����d�e�a�u�W�W�������]��G1�����9�2�6�d�m��3���>���F�UךU���:�&�4�!�6�����&����P9��N��1�����o�u�g�f�W�������R��V��!���d�3�8�e�m��3���>����v%��eN��Eʱ�"�!�u�|�m�}�G��I����W�=N��U���&�4�!�4��	��������\��c*��:���
�����m��������\�^�E��e�d�w�_�w�}��������C9��h��*���
�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����F�T�����u�%��
�#�����Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��n�u�u�6�9�)����	����@��Q��A��������4���Y����W	��C��\��u�e�e�e�f�m�G��Y����\��V ������&�c�3�:�h�Mύ�=����z%��r-��'���e�1�"�!�w�t�M���I����V��^�����u�:�&�4�#�<�(���
�ѓ�@��T��!�����
����_������\F��T��W��e�e�e�e�u�W�W�������]��G1��*���
�&�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����D��N�����!�;�u�%���ց�
����	F��s1��2������u�f�}�������	[�^�E��e�e�n�u�w�>�����ƭ�l5��D�*���
�u�u����>���<����N��
�����e�u�h�w�f�m�G��I����F�T�����u�%��
�#�l����H����`2��{!��6�����u�d�w�2����I����D��^�E��e�n�u�u�4�3����Y����\��h��G��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D��ۊ�u�u��
���(���-���F��@ ��U���o�u�d�n�w�}��������R��X ��*���g�f�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�e�e�d�l�}�WϽ�����GF��h�����#�g�c�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�d�g�f�W�������R��V�����
�#�g�b�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�f�l�L���YӅ��@��CN��*���&�
�#�g�n�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�F��Y����\��V �����:�&�
�#�e�e�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�G��B�����D��ʴ�
�:�&�
�!�o�6��*����|!��h8��!���}�d�1�"�#�}�^��Y����V��^�E��e�e�e�e�g�m�G��I��ƹF��X �����4�
�:�&��+�E��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������!�4�
�:�$�����M����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����4�!�4�
�8�.�(���K�Պ� %��N�&���������W��Y����G	�N�U��d�d�d�e�g�m�F��I����V��^�E��u�u�6�;�#�3�W�������l
��1��4����u�u����>���<����N��
�����e�u�h�w�g�l�F��I����V��^�D��d�d�d�w�]�}�W���
������T�����f�
�b�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�d�d�f�f�W�������R��V�����
�#�g�d�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�f�l�U�ԜY�Ư�]��Y�����;�!�9�m�g�g�$���5����l0��c!��]���:�;�:�e�w�`�U��I����]ǻN�����4�!�4�
�8�.�(���J���5��h"��<������}�e�9� ���Y���F�^�E��e�e�e�e�g�m�G���s���P	��C��U���6�;�!�9�f��G��Cӵ��l*��~-��0����}�a�1� �)�W���C���V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��Dߊ�a�e�o����0���/����aF�N�����u�|�o�u�f�m�F��I����V�=N��U���&�4�!�4��2����˹��\��c*��:���
�����}�������	[�_�D��w�_�u�u�8�.��������]��[�*��u�u��
���(���-���R��X����u�h�w�e�g�m�G��I����l�N�����;�u�%�6�9�)���&����	F��s1��2������u�f�}�������	[�^�E��e�e�e�e�l�}�WϽ�����GF��h�����#�`�a�e�m��3���>����v%��eN��Aʱ�"�!�u�|�m�}�G��H����V��^�����u�:�&�4�#�<�(���
����V��T��!�����
����_�������V�S��E��e�e�e�w�]�}�W���
������T�����d�
�u�u���8���&����|4�Y�����:�e�u�h�u�m�G��I����V��_�����u�:�&�4�#�<�(���
����^��rN�&���������W��Y����G	�N�U��e�e�e�e�f�l�F��[���F��Y�����%�6�;�!�;�n�(���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��I����9F������4�
��3�:�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��UךU���!�'�7�!�w�.�(�������\��C���ߊu�u�!�'�5�)�W���&����W��������3�8�o�$�:����
�Ģ�]�=N��U���;�9�4�
�>�����*����9��Z1�Oʆ�����]�}�W�������C9��P1����u�u����f�W���
����_F��1�����<�u�u����>���<����N��
�����e�n�u�u�$�:����&ù��C��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�<�;�;�-�G�������W9��h��U����
���l�}�Wϭ�����C9��v1��*���
�'�2�o���;���:���V�=N��U���;�9�%�d�:�%��������`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ�d�8�-�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���@��V��*ۊ�4�
�%�#�3�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�l��������W9��R	��U���
���u�j�z�P�ԜY�ƿ�T����*���<�1�<�
�>�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��1�����
�'�2�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�f�W���
����_F��1�����
�%�#�1�>�����Y����)��tUךU���<�;�9�%�e�����&����_��E��Oʆ�����m�}�G��Y����Z��[N��@���<�
�<�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�9��G��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�>�3�Ϯ�L����C9��S1��*���u�u��
���L���Yӕ��]��G1��7���
�9�
�'�0�g�$���5����\�^�����u�<�;�9�'�j�4���&����	F��s1��2������u�d�}�������9F������%�b��%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���@��V��*݊�
�%�#�1�>�����Y����)��tUךU���<�;�9�%�`���������V�=��*����u�h�r�p�W�W���������h��D���%�u�u����>���<����N��
�����e�n�u�u�$�:��������F��d:��9�������w�n�W������]ǻN�����9�4�
�<��.����&����U��N�&������_�w�}����Ӈ��@��U
��D���o�����W�W���������D�����
��&�b�1�0�A��*����|!��d��Uʦ�2�4�u�%�$�:����H���$��{+��N���u�&�2�4�w�-�������� W�,��9���n�u�u�&�0�<�W���������C1�*ۊ� �a�g�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����U5��z;��G���!�g�
�
�2��O���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N�����
�l�
�g�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������`9��b,�� ���f�'�2�a�a�g�$���5����l0��c!��]��1�"�!�u�~�W�W������� ��O#��!���!��9�<�;��@���&����CT�=��*����
����u�FϺ�����O��N�����4�u��-��	�8���4����C
��Y�����l�u�u����>���<����N��
�����e�n�u�u�$�:����	����l��F1��*���
�&�
�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�1��h�W���6����}]ǻN�����9�3�
���$��������_��1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������f*��x��8���<�9�
�a�%�:�C��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��&���1�
�0�8������5����E��h��*��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���
����@��d:�����3�8�l�o���;���:���F��P ��U���&�2�7�1�f�i�MϜ�6����l�N�����u�'�
�
���(���H�֓�C9��Y��U���
���n�w�}�����ƪ�l��R1������4�6���/����&¹��T9��N�&���������W��Y����G	�UךU���<�;�9�3��2��������~��d)�����<�d�g�'�0�h�F��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������
�0�8���?�$���
����lW��R	��D���u��
����2���+����W	��C��\�ߊu�u�<�;�;�:����I����l ��V�����!�'�u�u���8���B�����Y�����3�e�3�f�1��O߁�	����VF��d:��9����_�u�u�>�3�Ϲ�	����l ��h��D���4�
�0�1�w�}�#���6����9F������2�%�3�e�1�n����Aù��l��_��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���&����U��^�����-�g�o����0���/����aF�N�����u�|�_�u�w�4��������lV��h]�� ��e�<�
�0�6�m�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E��*ڊ�
�
� �d�g�<�(�������\��c*��:���
�����l��������l�N�����u�'�
�
���(���H�֓�C9��C��*���u��
����2���+������Y��E��u�u�&�2�6�}����&ù�� 9��h_�*���'�!�'�
�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����T��Q1�����3�
�m�
�'�/����&����`2��{!��6�����u�b�3�*����P���F��P ��U���
�
�
�
��(�F�������\��c*��:���n�u�u�&�0�<�W���
����@��d:��ӊ�&�
�u�u���8���B�����Y�����<�
�1�
�n�}�W���5����9F������2�%�3�e�1�i����AĹ��l��E��U���
���n�w�}�����ƫ�C9��1��A���
�m�
�%�3�3�W���-����t/��=N��U���;�9�2�%�1�m��������9��h���������W�W���������h��*���
� �d�b�6�����Y�Ɵ�w9��p'�����u�<�;�9�0�-�����ғ�F9�� 1��*���'�0�!�e�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��h^��*ފ� �d�b�<��8����J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�
�
�
��(�F�������V��Y��U����
�����#���Q����\��XN�N���u�&�2�4�w�/�(���&����U��Y�����0�6�;�
�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����T��Q1�����3�
�m�
�'�/����&����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʲ�%�3�e�3�c�;�(��&����V��Y1�Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-�����ғ�F9�� 1��*��� �;�g�o���;���:����g)��]����!�u�|�_�w�}����Ӂ��l ��h��*���d�b�4�
�2�(���Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
�
�
�
�"�l�@���&����A��T��!�����
����_������\F��d��Uʦ�2�4�u�'���(���&����Q��G1�����
�u�u����>���<����N��
�����e�n�u�u�$�:��������9��1��*��
�%�6�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�&�&��(���H����lW��N��1�����_�u�w�4��������T9��S1�G������]�}�W�������A��h^��*ي� �d�e�4��)����	����A��R	��U���
���u�j�z�P�ԜY�ƿ�T��	��*���
�
�
� �f�j��������R��C��*���u�u��
���W��^����F�D�����'�
� �d�b�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����l�
�d�o���;���:����g)��]����!�u�|�_�w�}����Ӈ��@��T��*���&�g�3�8�f�g�$���5����l�N�����u�%�&�2�5�9�E��CӤ��#��d��Uʦ�2�4�u�%�$�:����&����GS��D��U����
���l�}�Wϭ�����R��^	�����`�u�u����L���Yӕ��]��P�����l�
�e�o���;���:����g)��]����!�u�|�_�w�}����Ӂ��l ��W�����u��
����2���+������Y��E��u�u�&�2�6�}�$���,����F��B�����d�
� �g�d�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��Q=��8���,� �
� �#�-���&����U��N�&���������W��Y����G	�UךU���<�;�9�3���;�������_��[��A���
�e�
�e�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������`9��b"��:����9�<�9��i����I˹��\��c*��:���
�����l��������l�N�����u�
�4�g�$�;�(��&���5��h"��<������}�f�9� ���Y����F�D�����:�
�
� �e�i����Y����)��t1��6���u�b�1�"�#�}�^�ԜY�ƿ�T����*���
� �g�a�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1�����g�
� �g�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��*���
� �g�m�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��*��� �g�e�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����G�� V��*���
� �g�m�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��D���3�
�m�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��*��� �g�c�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V��h��*���4�!�6�&��(�E���	����`2��{!��6�����u�d�w�2����I��ƹF��^	��ʦ�9�!�%�<�1��@݁�J����g"��x)��*�����}�a�3�*����P���F��P ��U���0� �!�&�1��G߁�J����g"��x)��*�����}�b�3�*����P���F��P ��U���-� ��;�"��G���&����e9��Q��EҊ�g�o�����4���:����W��S�����|�_�u�u�>�3�Ϫ�	�Փ�l ��_�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)�������� T��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�a�
� �d�m����Y����)��t1��6���u�b�1�"�#�}�^�ԜY�ƿ�T����*���3�
�a�
�f�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��\�� ��g�%�u�u���8���&����|4� N�����u�|�_�u�w�4����	����9��^1��*��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������l��B1�E���u�u��
���(���-��� V��X����n�u�u�&�0�<�W�������lW��Q��CҊ�`�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�&����gT��B��E���
�%�,�0�1��N݁�J����g"��x)��*�����}�a�3�*����P���F��P ��U���
�8�c�<�1��Oہ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�
�
�"�n�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����8�m�<�3��d�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*����g��!�e����I����	F��s1��2������u�d�}�������9F������2�%�3�
�n����*����|!��d��Uʦ�2�4�u�%�$�:����&����GP��D��U����
���l�}�Wϭ�����R��^	�����a�u�u����L���Yӕ��]��P�����l�
�0�o���;���:���F��P ��U����
�&�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƭ�l��h��*���o�����W�W���������D�����g�a�o����9�ԜY�ƿ�T�������7�1�`�u�w��;���B�����Y�����<�
�1�
�d�g�5���<����F�D�����%�&�2�7�3�j�W���6����}]ǻN�����9�4�
�<��9�(��CӤ��#��dךU���:�%�;�;�w��B���8����l ��'��U���%�'�u�_�w�}�W���	����\��yN��1�����_�u�w�}�W������/��d:��9����_�u�u�w�}�������/��d:��9����_�u�u�w�}��������|3��d:��9����_�u�u�w�}��������|3��d:��9����_�u�u�w�}�������)��=��*����n�u�u�w�}��������F��~ ��!�����
����_������\F��d��U���u�<�
�4��}�W���*����|!��h8��!���}�d�1�"�#�}�^�ԜY���F��h����o��u����>���<����N��
�����e�n�u�u�w�}��������lV�!��U���
���
��	�%���Hӂ��]��G�U���u�u�4�
�2�(���Cө��5��h"��<������}�f�9� ���Y����F�N�����0� �;�g�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y���R��R����o������0���/����aF�
�����e�n�u�u�w�}��������}F��s1��2���|�_�u�u�9�}��������9lǻN�����;�;�u��b�j�6���I����/��N�����u�_�u�u�w�}��������}F��s1��2���_�u�u�u�w�-����Cӯ��`2��{!��6�ߊu�u�u�u�'�.����Cӯ��`2��{!��6�ߊu�u�u�u�'�9����Y����`2��{!��6�ߊu�u�u�u�'�4����Y����`2��{!��6�ߊu�u�u�u�'�/����Cө��5��h"��<��u�u�u�u�>���������\��yN��1��������}�D�������V�=N��U���u�;��'�8��W���7ӵ��l*��~-��0����}�d�1� �)�W���s���F�^ �����0�!�d�o��}�#���6����e#��x<��F���:�;�:�e�l�}�W���Yӏ��d��T��*���u������4���:����U��S�����|�_�u�u�w�}��������F��x;��&���������W��Y����G	�UךU���u�u�%�'�#�/�(���Y����`2��{!��6�����u�f�w�2����I��ƹF�N�����!�'�
�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����C9��C��*���u� �u����>���<����N��
�����e�n�u�u�w�}��������lR�!��U���
���
��	�%���Hӂ��]��G�U���u�u�4�
�2�(���Cө��5��h"��<������}�f�9� ���Y����F�N�����0�o��u���8���Y��ƹF��Y
�����;�;�n�_�w�}����������/��4���e�3� �
�e�.�Dݰ�&�ԓ�l ��[1��ʜ�_�u�u�0�2�4�W�ԜY���F��T��;����n�u�u�w�}�9���*����\��y:��0��u�u�u�u�3�3�(���-����z(��p+�����u�u�u�<�f�
�3���Cӯ��v!��d��U���u�1� �
��	�W���7����aF�=N��U���!�}�u�u�w�}����Cӯ��`2��{!��6�ߊu�u�u�u�2�8�W���7ӵ��l*��~-�U���u�u�1�;�w�}�9ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y���W��T��;ʆ�������8���J�ƨ�D��^����u�u�u�0�m��W���&����p]ǻN��U���:�!�o����3���>����v%��eN��Dʱ�"�!�u�|�~�W�W����Ư�^��R ���ߊu�u�:�%�9�3�W���L�щ�p ��h����;�
�g�&�d��(���&����z5ǻN�����<�u�_�u�w�}�W���Cӯ��v!��d��U���u������Mϗ�-����l�N��Uʱ�;�
���w�}�9���<��ƹF�N��������o��	�0���s���F�S��*����u�u����W��Y����\��d��U���u�1�;�u�w��$���5����l0��c!��]��1�"�!�u�~�W�W���Y�ƨ�]W�'��&���������W��Y����G	�UךU���u�u�:�!�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�^�ԜY�Ʃ�WF��Z�����_�_�7�2�9�}�WϹ�	����l ��h��D��o�6�8�:�2�)���8ģ��U9��Q1�U���%�'�u�4�w�W�W���Y�ƭ�l��S����9�y�u�u�w�}����
�����E�����u�u�u�%�$�<���Y����U9��Q1�����m�
�%�&�6�)�}���Y���R��X ��H���'�
�
�
�����I����W	��d��U���u�4�
�1�2�`�W���&����U9��Q��Mڊ�%�<�9�y�w�}�W�������R��
P�����
�
�
�
�"�l�G���&����JJǻN��U���;�4�%�4�f�`�W���&����U9��Q��Mڊ�;�4�%�4�f�W�W���Y�ƥ�l��h\��Kʲ�%�3�e�3�d�;�(��&����R��d��U���u�<�
�0�6�m�J�������9��1��*��
�;�7�!��q�W���Y����C9��C��*���k�2�%�3�g�;�D���&����R��R����_�u�u�u�w�-��������X��E��*ڊ�
�
� �d�g�<�(�������l�N��Uʴ�
�0� �;�e�`�W���&����U9��Q��Mڊ�%�'�!�'��q�W���Y����C9��C��*���k�2�%�3�g�;�D���&����R��R����_�u�u�u�w�-����GӁ��l ��h��*���d�e�4�
�2�f�}���Y����U9��Q1�����m�u�u�:�'�3����<�Ӎ�v'��h^��*�ߊu�u�:�!�:�-�_���Y�����T��H���%�6�>�_�w�}�W���	����[�V�����u�u�u�u�6�����Y����A��h^��*ފ� �d�b�4��)���Y���F��G1�����k�2�%�3�g�;�C���&����R��X �����u�u�u�%�>�1�W�������lV��hZ�� ��b�4�
�1�2�W�W���Y�ƭ�l��S��Kʲ�%�3�e�3�c�;�(��&����V��d��U���u�<�
�%�%�8���D�ƫ�C9��1��A���
�m�
�;��8����&��ƹF�N�����'�:�
�u�i�:����I����l ��V�����0�<�1�f�]�}�W���Y����C��R ��D��u�'�
�
���(���H�ѓ�]9��R�����y�u�u�u�w�4�(�������lT�	N�����e�3�a�3��e�(���.����V��BךU���u�u�%�'�#�/�(���GӁ��l ��h��*���d�b�4�
�2�(���s���F�V�����;�d�h�u�%��(߁�&ǹ��lW��h�����'�
�y�u�w�}�WϿ�&����A��S����3�e�3�a�1��O؁�	����F��BךU���u�u�%�'�#�/�(���GӁ��l ��h��*���d�b�4�
�2�(���s���F�V�����;�a�h�u�%��(߁�&ǹ��lW��h�����'�
�y�u�w�}�WϿ�&����A��S����3�e�3�a�1��O؁�	����F��BךU���u�u�%�6�w�c�����֓�lR��B1�B���
�0�n�_�w�}�(߁�
������\��*���f�3�9�
�$��F���Y����\��CN��Eߔ���
�
�$�?�Dݰ�&�Ԣ�lU��1�����&�_�u�u�2�8�������F�N��<���k�d�_�u�w�}�W���&����vF�]�U���u�u�1�;���#���G����9F�N��U���d����j�}�E�ԜY���F��B��<���u�k�f�|�w�}����Y����l�N��Uʶ�>�h�u�%�4�6�}���Y���A��CN��U���'�!�_�u�w�}�W���I���T��Q��Lߊ�e�_�u�u�w�}���D�ƫ�C9��h_�*��_�u�u�u�w�8�J�������lW��h�����u�u�u�:�#�`�W���&����
S��G����u�
�
�&�5�n����K����9��Q��*���
�d�u�u�8�-����Y����rQ��t��*���7�f�;�
�e�.�D݁�&����l��=N��U���0�<�u�4�w�W�W���Y�ƅ�[�BךU���u�u� �
���W���J���F�N��ڊ���u�k�d�q�W���Y����Z��`'��=��u�g�_�u�w�}�W�������g.�	N�\���u�%�'�u�6�}�}���Y���P
��
P�����>�_�u�u�w�}����Y����C9��CBךU���u�u�<�e�j�}��������l��=N��U���u�<�d�h�w�/�(���H�ߓ�JǻN��U���0�h�u�'��(�F�����ƹF�N�����h�u�'�
�"�l�N���P��ƹF��h^�����f�;�
�g�$�n�(ށ�����C9��N����:�0�!�8�g��2���&ù��F
�� ��Fػ�
�g�d�8�/�9����YӁ��V����U�ߊu�u�u�u��`�W��Y���F��b#��!���u�k�d�_�w�}�W����֓�z"��S�F���u�u�u�u�3�3�(���-���U��=N��U���u�:�!����J���K���F��E�����_�u�u�u�w�4�G��Y����~3��N!��*���!�%�,�d��(�E���	��ƹF�N����h�u��-��	�8���4����C
��Y�� ��f�%�y�u�w�}�WϺ���� ��O#��!���!��9�<�;��@���&����CT�=d��Uʳ�e�3� �
�e�.�Dݰ�&�ԓ�l��h
��*��u�u�:�%�9�3�W���L�щ�p ��h����;�
�g�&�d��(���&����F�P�����8�%�}�u�w�}�Wϗ�Y���l�N��Uʛ�����j�}�[���Y�����1��1���h�u�g�_�w�}�W����ד�z"��S�F���u�u�u�u�3�(�(���-���U��=N��U���!�8�%�}�w�}�W�������X��d1�� ����!��9�>�1�(�������9��d��U���u�1�;�u�i�;�(���5����G9��[�����a�3�
�e��l�}���Y���W	��S������,� ��(���� ����U��V��G��_�_�_�u�w�p��������]��C��U´�
��3�8�w�;����
������_��[���_�u�u�%������
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��h-�����i�u�%���)�(���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�V�N��U���u�u�u�u�w�}����*����Z�V��&���8�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��E��*ڊ�
�
� �d�g�<�(�������l��E�����&�<�;�%�8�8����T�����h��*���
� �d�e�6�����&����G��h��*���<�;�%�:�w�}����
�έ�l��d��Uʷ�2�;�u�u�w�}��������XA��R �����4�
�9�u�w�z�P�����ƹF�N��U���3�}�%�'�#�`�P���Y����9F�N��U���u�u�u�'���(���&����V��G1�����4�
�!�'��8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�n�;���P�Ƹ�V�N��U���u�u�u�u�w�}�����֓�lU��B1�E���
�!�'�
�'�.�������F��h�����:�<�
�n�w�}�W���Y���F��[��U���%�6�;�!�;�:���DӁ��l ��h��*���d�e�4�
�2�9�^������F�N��U���u�u�u�u�0�-�����Փ�F9��1��*���'�
�%�&�6�)����E�ƭ�l��D�����
�n�u�u�w�}�W���Y����]��QU��U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K�P�����3�a�3�
�o���������C9��V�����4�&�2�u�%�>���T���F��G1��E���a�3�
�m��-��������@��C1�����&�2�
�'�4�g��������C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�}�F�������F�N��U���<�u�4�
�$�}�W��PӒ��]l�N��U���u�u�u�2�'�;�G���M����^��V�����
�%�&�4�#�/���Y����\��h�����n�u�u�u�w�}�Wϻ�
���F�N��U���u�<�u�}�6�����&����P9��
N��*���u�;�u�4��2��������F�V�����&�$��
�#�m����@�ƭ�WF��CF�����;�!�9�2�4�m�JϹ�	����l ��h��D���4�
�:�0�~�t����Y���F�N��U���u�u�u�'���(���&����Q��G1�����4�
�!�'��8�W������]��[����_�u�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����&ù��9��h_�*���'�4�,�|�#�8�W���Y���F�N��U���u�'�
�
���(���H�ѓ�C9��V�����!�'�
�0�w�`��������_	��T1����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l'��G1�����0�u�&�<�9�-����
���9F���*���%�#�1�%�2���������PF��G�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�I�����_�u�u�u�w�}�W���Q����@�I�\ʡ�0�_�u�u�w�}�W���Y�Ƽ�9��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W�������C9��P1����a�u�=�;�]�}�W���Y���F�N��U���%�e��4��1�(������R��X ��*���<�
�n�u�w�}�W���Y���F������4�
�<�
�3��B������F�N��U���u�u�u�u�w�}����8����E
��G��U��%�e��4��1�L���Y���F�N��U���u�;�u�3�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���
�
�'�2�6�.��������@H�d��Uʥ�e��%�0��.����	����	F��X��´�
�9�|�u�w�?����Y���F��QN�����>�0�0�!�6�9�������A��N���ߊu�u�u�u�w�}����	����[�I�����_�u�u�u�w�}�W���Y����r9��R	��Hʴ�
�:�&�
�!�o�G�ԜY���F�N���ߊu�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�
�������ƭ�WF��CF�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�6�9�_�������l
��^��U���%�&�4�!�~�t�W������F�N��U���u�u�u�%�g�����Y����lV��d��U���u�u�u�u�w�8�Ϸ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�Z���&¹��K9��h��*���2�4�&�2�w�/����W���F�G1�����4�
�9�
�%�:��������\������}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�_��U���;�u�u�u�w�}�WϷ�Yۇ��A��
N��R���=�;�u�u�w�}�W���Y����lW��V�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƥ�N��h��*���
�f�|�!�2�}�W���Y���F�N��U���u�u�
�
�6���������TF������!�9�2�6�g�W�W���Y���F�N��Uʰ�&�3�}�%�$�:����L����[��=N��U���u�u�u�u�w�}�W���Y����^��V�����'�2�i�u������	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�f�0�����ƭ�@�������{�x�_�u�w��(���&����l��^	�����u�u�'�6�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�r�r�u�?�3�W���Y���F��QN�����!�h�r�r�w�5����Y���F�N��U���
�4�
�'�0�a�W�������l
��1����u�u�u�u�w�1����Y���F�N��U���}�}�%�6�9�)���������T�����;�!�}�4��2��������F�V�����&�$��
�#�����PӇ��N��h�����:�<�
�u�w�-�������R�������!�9�2�6�f�`��������C9��SG��U���;�_�u�u�w�}�W���Y���F��1�����0�u�h�%�f�0��ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
�2�4����&����C�������%�:�0�&�w�p�W���	�ԓ�V��S1��*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�K����Z	��V�����'�2�i�u�'�>��������lV��N��U���u�u�0�&�]�}�W���Y���F�^��]���6�;�!�9�0�>�F������O��_��U���u�u�u�u�w�}�W�������C9��P1����a�u�=�;�]�}�W���Y���F�N��U���%�g��'�8���������TF������!�9�2�6�g�W�W���Y���F�N��Uʰ�&�3�}�%�$�:����O����[��=N��U���u�u�u�u�w�}�W���Y����c��X
�����1�%�0�u�j�-�E�������R��[
�U���u�u�u�u�w�}�W�������U]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p����)����W9��R	�����;�%�:�0�$�}�Z���YӖ��l6��^�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��(�������A��S�����;�!�9�f��f�W���Y���F��[��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}�������R��X ��*���<�
�u�u�'�.��������l��h��*���4�1�}�%�4�3��������[��G1�����|�u�;�u�6�����&����P9��
N��G���'�:�
�%�!�9�^������F�N��U���u�u�u�u�'�o�'�������V�
N��G���'�:�n�u�w�}�W���Y�������U���u�u�u�u�w�8�Ϸ�B���F���U���_�u�u�;�w�/����B��ƹF�N��@���4�
�9�
�%�:�����Ƽ�\��D@��X���u�%�`��6���������@��Y1�����u�'�6�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���r�r�u�=�9�}�W���Y����������h�r�r�u�?�3�W���Y���F�N��*ߊ�
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W������F�N��U���u�3�}�4��2��������F�V�����!�0�_�u�w�}�W���Y���F�^�����<�
�1�
�d�t����Y���F�N��U���u�u�u�u�w��(���	����l��PN�U���6�;�!�9�0�>�G�ԜY���F�N��U���u�0�&�3��-��������O��_�����u�u�u�u�w�}�W���Y���C9��u1��*���
�'�2�i�w��(���	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�b�����Y����T��E�����x�_�u�u���(�������Z��G��U���'�6�&�}�'�>��ԜY�Ʈ�T��N��U���<�u�4�
�;�z����Y����R��[��U��r�u�=�;�w�}�W���Y����UF��G1����r�r�u�=�9�}�W���Y���F���*���'�2�i�u�'�>��������]ǻN��U���u�u�9�0�w�}�W���Y���F��QN��]���6�;�!�9�0�>�F������F��SN�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^�������C9��Y�����6�d�h�%�b����������YNךU���u�u�u�u�w�}�W���&ƹ��C��R������_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��hY��*���#�1�%�0�w�.����	����@�CךU���
�
�
�%�!�9����&����T��E��Oʥ�:�0�&�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��U��|�!�0�_�w�}�W���Y�ƥ�N��h��U���d�|�!�0�]�}�W���Y���F�G1��6���
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y����������7�1�g�a�w�5��ԜY���F�N��U���u�u�u�%�`���������V�
N��*���&�
�:�<��f�W���Y���F�N��U���9�<�u�4��4�(���&���G��d��U���u�u�u�u�w�}�W���YӖ��l%��G1�����0�u�h�%�`�������ƹF�N��U���u�u�u�u�9�}��ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�
��/�Ͽ�
����C��R��U���u�u�%�b��-����
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F�� 1�����u�h�4�
�8�.�(���K����F�N��U���0�&�_�u�w�}�W���Y���Z �F��*���&�
�:�<��}�W�������]��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
��-����P�Ƹ�V�N��U���u�u�u�u�w�}����:����TF���*��u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���R��P �����&�{�x�_�w�}����
����C9��\GךU���0�<�_�u�w�}�W���Q����_��A��U���u�%�6�>�j�z�P�����ƹF�N��U���3�}�}�%�4�3��������[��G1��\ʴ�1�}�%�6�9�)���������D�����
��&�d��.�(�������\�V�����
�:�<�
�w�}����&ù�� 9��h_�*���1�;�|�|�w�5����Y���F�N��U���;�1�
�0�:��:���*����A��h_��*���
�e�u�h�0�-�����Փ�F9��1��*��� �;�d�_�w�}�W���Y���F��h �����'�
��4�4��(�������9��P1�D��u�'�
�
���(���H�֓�C9��C��*��u�u�u�u�w�}�W�������W��R��&���7���&�4�4�F�������Z�P�����3�f�3�
�o���������]ǻN��U���u�u�u�u��3��������e+��T=��*���#�
�
�0��l�W������lV��h]�� ��e�4�
�0�"�3�D�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�<����Y����V��C�U���%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z �F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h_��U���6�|�4�1�9�)��������W9��G��U���;�u�u�u�w�}�W���YӀ��K+��c\�� ���e�d�'�2�c�l�K���*����2��x��Gڊ�
� �a�g�'�f�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠu�u�x�u�$�4�Ϯ�����F�=N��U���6�&�u�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��R��u�=�;�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1����|�u�=�;�w�}�W���Y���F��d1�� ����!��9�>�1�(�������
P�
N��*����,� �
�"�)����Hǹ��lT��h����u�u�u�u�w�}�W�������J)��h#�����,�d�
�0��d�W������f*��x��8���<�9�
�b�1��G܁�K���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���6�&�n�_�w�}�ZϿ�
����C��R��U���u�u�%�:�2�.�_������F�U�����u�u�u�<�w�<�(���^����GF��SN��*���u�u�d�|�#�8�}���Y���F�^��]´�
�:�&�
�8�4�(���Y����VO��Y
�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�~�)��ԜY���F�N��Uʳ�
����#�o�(���&����[��E�� ��l�%�n�u�w�}�W���YӃ����=N��U���u�;�u�3�]�}�W���Y����V��=d��U���u�&�<�;�'�2����Y��ƹF��E�����4�
�9�|�w�}�������F���]���6�>�0�0�#�<�Ͽ�&����F�G�����u�u�u�u�w�}����Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��h]��U���}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�^�����ƹF�N��U���u�u�0�
�f�}�JϹ�	����_��G\�U���u�u�u�u�2�9���Y���F��Y
���ߊu�u�;�u�%�>���s���K��_�����&�4�0�}�'��(���PӉ��G��D��ʸ�6�<�0�u�z�}�WϿ�&����@��D�����:�u�u�'�4�.�Wǿ�&����@�V�����%�&�2�7�3�l�F�������9��1��*��
�%�1�;�{�:����I����l ��V�����:�0�_�u�w�8��ԜY���F��D�����
�&�u�&�w�}�W���Y����[��V��!���d�3�8�e�j�}�W���Y���F�N�����}�%�6�;�#�1����H����C9��N��ʻ�!�4�
�<��9�(��P����[��N��U���u�u�u�u�w�}����*����Z�V��!���g�3�8�d�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:��؊�&�
�u�k�]�}�W���Y���F�V��&���8�i�u�%���܁�
����9F�N��U���u�=�;�4��	��������[�=N��U���u�u�u�u�w�-�9���
�����d:��ފ�&�
�n�u�w�}�W���Yӑ��]F��h=�����3�8�f�h�w�}�W���Y���F���;���&�u�h�4��	��������l�N��U���u�"�0�u�'��(���&����F�d��U���u�u�u�u�w�<�(������F��h=�����3�8�`�_�w�}�W���Y�ƻ�V��G1��*���
�&�
�u�i�W�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�=�;�6��#���N����lP�	NךU���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y����[��V��!���m�3�8�b�j�}�W���Y���F�N�����
�&�u�h�6��#���@����l^��N��U���u�u�"�0�w�-�$���ʹ��^9��
P��U���u�u�u�u�w�}����*����Z�V��!���d�
�&�
�l�}�W���Y�����YN��*���&�d�
�&��}�I�ԜY���F�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�:�}�4��2��������F�P�����3�f�3�
�o��������F��R ךU���u�u�u�u�w�}�W���	����U��S�����
�!�d�3�:�l�L���Y���F�N��U���0�u�u�u�w�}�W���Y�����y=�����h�4�
��$�l�(���&��ƹF�N��U���u�u�;�u�1�W�W���Y���F��R �����
�!�d�3�:�l�W���s���F�N��U���<�u�}�4��2��������F�V�����;�u�:�}�6�����&����P9��
N�����e�3�a�3��e�(�������O�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���0�u�u�u�w�}�W���Y�����y=�����h�4�
��$�l�(���&����F�N��U���u�u�0�1�>�f�W���Y���F��_�����'�u�k�u�w�}�W���Y���F��G1��*���u�h�w����/���[���F�N��ʶ�&�n�u�u�2�9��������9F�C����:�0�4�&�0�}����
���l�N��*���0�4�&�2��/���	����@��G1��Yʲ�%�3�e�3�c�;�(��&����\�������6�0�
��$�l�(���&���F�U�����u�u�u�<�w�u��������_	��T1�Hʴ�
�0�u�;�w�<�(���
����T��N�����<�
�&�$����������O��Y
�����4�
�:�&��2����Y�ƫ�C9��1��A���
�m�
�%�3�3�^���Y����l�N��U���u�4�
�:�2�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���<�9�u�&�>�3�������KǻN�����9�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��GךU���0�<�_�u�w�}�W���Qۈ��N��h�����:�<�
�u�w�-��������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�|�!�2�}�W���Y���F��G1�����h�4�
�:�$�����&��ƹF�N�����_�u�u�u�w�}�W�������[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���T�ƭ�l��S�����;�%�:�0�$�}�Z���YӇ��A��N1�����
�'�6�o�'�2��������F��G1��E���a�3�
�m��-����UӇ��@��T��*���&�d�
�&��m�}���Y����]l�N��Uʼ�u�}�4�
�8�.�(�������F��h��U���u�4�
�:�$�����&���R��^	������
�!�d�1�0�F�������\�V�����
�:�<�
�w�}����&ù��9��h_�*���1�;�|�|�w�5��ԜY���F�N��*���1�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����V��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����1�d�`�4�$�:�W�������K��N�����<�
�1�
�g���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����I���N��h�����#�
�u�u�'��(���Q�ƨ�D��]��N���u�0�1�%�8�8��Զs���K��G1�����1�d�a�4�$�:�W�������K��N�����<�
�1�
�f���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����H���N��h�����#�
�u�u�'��(���Q�ƨ�D��X��N���u�0�1�%�8�8��Զs���K��G1�����1�d�d�4�$�:�W�������K��N�����<�
�1�
�d���������PF��G�����4�
�!�'�{�-�G�������W9��h��Yʥ�d�8�-�4��1�(���
���C9��g�����%�#�1�<��4�[Ϯ�L����C9��S1��*���y�%�b��6���������l�N�����u�u�u�u�w�}�W�������T9��S1�D��u�}�
�
��-��������TF�V�����
�:�<�
�~�2�WǮ�L����C9��S1��*���u�u�%�6�9�)�������\�G1��%���:�
�%�#�3�4�(���Y�ƭ�l��D�����
�|�:�u�'�l��������W9��h��U���%�6�;�!�;�:���Y���C9��v1��*���
�;�&�2�j�<�(���
����T��G�����%�&�4�!�j�<�(���
����T��G����u�;�u�'�4�.�L�ԶY���F��h��*���
�`�u�&�>�3�������KǻN�����2�7�1�d�e�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���K�����T�����d�d�h�4������Nӂ��]�� G����u�;�u�'�4�.�L�ԶY���F��h��*���
�c�u�&�>�3�������KǻN�����2�7�1�d�c�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���M�����T�����d�d�h�4������@ӂ��]��G����u�;�u�'�4�.�L�ԶY���F��h��*���
�l�u�&�>�3�������KǻN�����2�7�1�d�b�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���L�����T�����d�d�h�4������Aӂ��]��G����u�;�u�'�4�.�L�ԶY���F��h��*���
�g�u�&�>�3�������KǻN�����2�7�1�g�e�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���K�����T�����d�d�h�4������H�ƨ�D��_�\�ߊu�u�;�u�%�>���s���K�V�����1�
�f�u�$�4�Ϯ�����F�=N��U���&�2�7�1�e�i��������\������}�'�
�
���(���H�ѓ�C9��Y����<�
�&�$����������OǻN�����_�u�u�u�w�}�W���Y����Z��S
��F���h�}�4�
�8�.�(�������F��h��*���$��
�!�f�;���PӇ����F��*���&�
�:�<��}�W���&����U9��Q��M݊�%�1�;�|�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����M�ƭ�@�������{�x�_�u�w�-��������^��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��A���h�}�%�6�9�)����H����C9��h��]���:�;�:�d�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����L�ƭ�@�������{�x�_�u�w�-��������S��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��@���h�}�%�6�9�)����H����C9��h��]���:�;�:�a�~�W�W����Ƽ�\��DUװ���u�x�4�
�>�����NӇ��Z��G�����u�x�u�u�6���������l��^	�����u�u�'�6�$�u����&����9F����ߊu�u�u�u�w�}�W���	����l��h\�I���4�
��3�:�m��������[��G1�����9�d�d�n�w�}����	����@��=d��U���u�%�&�2�5�9�C������]F��X�����x�u�u�4��4�(���&����R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��Z�I���4�
�:�&��+�(���Y����`9��ZF����!�u�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�C���
������T��[���_�u�u�%�$�:����Mƹ��@��h����%�:�0�&�6�����UӇ��@��T��*���&�d�3�8�g�}�(߁�&����_�N�����;�u�u�u�w�}�W���YӇ��@��U
��A���h�}�4�
�8�.�(�������F��1�����9�|�4�1�9�)�_ǿ�&����G9��P��D��4�
�<�
�$�,�$���¹��^9����U´�
�:�&�
�8�4�(���Y����G��G��N���u�0�1�%�8�8��Զs���K��G1�����1�`�u�&�>�3�������KǻN�����2�7�1�`��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����u�
�
�4��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����R�
N�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u������	����O��N�����%�:�0�&�]�W�W���TӇ��@��U
��C���&�<�;�%�8�8����T�����D�����c�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*؊�0�<�1�4��1�^���Yӄ��ZǻN��U���u�u�u�u�'�.��������[�Y��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�<����	����@��X	��*���u�%�&�4�#�t�W���Yۇ��P	��C1�����d�h�%�g��/����	����O��N�����%�:�0�&�]�W�W���TӇ��@��U
��B���&�<�;�%�8�8����T�����D�����b�
�&�<�9�-����Y����V��V�����y�4�
�<��.����&����U��B��*ߊ�
�%�#�1�]�}�W������F�N��U���u�4�
�<��9�(��E����\������!�9�2�6�f�`��������V��c1��D���8�e�u�;�w�<�(���
����T��N�����!�'�|�|�6�9�_�������l
��^��U���
�
�
�%�!�9�^�ԜY�Ʃ�WF��X���ߠ_�u�u�x�6�����������^	�����0�&�u�x�w�}��������W9��h�����%�:�u�u�%�>����	����A�V�����&�$��
�#�����UӖ��l%��G1���ߊu�u�0�<�]�}�W���Y���F�V�����1�
�l�i�w�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\ʴ�1�}�%�6�9�)���������h-�����1�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�&�&��(���I����l_��D��ʥ�:�0�&�u�z�}�WϿ�&����P��h=����
�&�
�
�$�4��������C��R�����<�
�1�
�a�t�W�������9F�N��U���}�%�&�2�5�9�F��Y����l�N��U���u�4�
�<��.����&����l ��hW��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��C_�����l�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�<�
�$�,�$����ד�@��N�����u�'�6�&�y�p�}���Y����Z��D��&���!�d�3�8�f���������PF��G�����4�
�<�
�3��E���Y����V��=N��U���u�3�}�%�$�:����K���G��d��U���u�u�u�4��4�(�������@��h��*��i�u�%�6�9�)��������F�N�����u�u�u�u�w�}�WϿ�&����P��h=����
�&�
�e�k�}��������\��h^�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�4��4�(�������@��Q��Eʴ�&�2�u�'�4�.�Y��s���R��^	������
�!�
�$��(�������A	��N�����&�4�
�<��9�(��s���Q��Yd��U���u�<�u�4��4�(���&���G��d��U���u�u�u�4��4�(�������@��Q��E��u�%�6�;�#�1����H���F�N�����u�u�u�u�w�}��������V��c1��D���8�e�i�u�'�>��������lV��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�4�
�<��.����&����U��N�����u�'�6�&�y�p�}���Y����Z��D��&���!�
�&�
��.����	����	F��X��´�
�<�
�1��i�^���Yӄ��ZǻN��U���3�}�%�&�0�?���A�Ƹ�V�N��U���u�u�4�
�>�����*����9��Z1�I���%�6�;�!�;�:���s���F�R��U���u�u�u�u�w�<�(���&����l5��D�����d�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]Ǒ=N��U���4�
�<�
�$�,�$���ǹ��^9��V�����'�6�&�{�z�W�W���	����l��F1��*���
�&�
�
�$�4��������C��R�����<�
�1�
�g�t�W�������9F�N��U���}�%�&�2�5�9�F��Y����l�N��U���u�4�
�<��.����&����U��N�U���6�;�!�9�0�>�F�ԜY���F��D��U���u�u�u�u�6�����
����g9��1����i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�&�&��(���&����F��D��U���6�&�{�x�]�}�W���
����@��d:��ߊ�&�
�
�&�>�3����Y�Ƽ�\��DF��*���
�1�
�`�~�}�Wϼ���ƹF�N�����%�&�2�7�3�o�B������F�N��U���4�
�<�
�$�,�$���ƹ��^9��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�4��4�(�������@��Q��A��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���ف�
����R��P �����&�{�x�_�w�}��������B9��h��*���
�
�&�<�9�-����Y����V��V�����1�
�a�|�w�}�������F���]���&�2�7�1�c�j�W������F�N��Uʴ�
�<�
�&�&��(���&����F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�4�
�>�����*����9��Z1�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���
�&�$���)�(���&�ƭ�@�������{�x�_�u�w�-��������`2��CY�����
�&�<�;�'�2�W�������@N��h��*���
�d�|�u�w�?����Y���F��QN�����2�7�1�d�c�}����s���F�N�����<�
�&�$���؁�
����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����U��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�V�����&�$��
�#�����Y����T��E�����x�_�u�u�'�.��������l��h��*݊�&�<�;�%�8�}�W�������R��^	�����`�|�u�u�5�:����Y����������7�1�d�g�w�5��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�d�_�w�}�W������F�N��U���4�
�<�
�$�,�$���˹��^9��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h��*���$��
�!��.�(���
������T��[���_�u�u�%�$�:����&����G_��D��*���<�;�%�:�w�}����
�έ�l��h��*��|�u�u�7�0�3�W���Y����UF��G1�����1�d�`�u�?�3�}���Y���F�V�����&�$��
�#�����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�<�
�&�&��(���&����F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y����~3�� ����
�
� �a�e�-�W��s���F�Q=��8���g��!�g��(�D���	�ƻ�V�D�����
�
� �f�a�-�_���D����F��D��U���u�u�%�e��4�(���B��� ��O#��!ػ� �
�e�3��e�(��E�Ƽ�a��[��M���
�c�
�`�]�}�W���������C1�*���0�%��d�1��Gׁ�K���@��[�����6�:�}�;�>�3�Ǯ�+����G9��Q��Eڊ�f�u�u�;�>�3�ǿ�&����G9��V��\��u�u�3�
���E�������Z��G:�����
�l�
�f�k�}�W���Y����V��h��*���4�!�6�&��(�E���	�ƻ�V�D�����
�
� �g�a�-�_���D����F��D��U���u�u�&�9�#�-����&����CU��N�������,� ��(���� ����U��V��E��u��-� �.�(�(�������P��N�������,� ��(���� ����U��V��D��u�%�6�;�#�1�D݁�<����r$��N�������,� ��(���� ����U��]��E��u�0�
�d�l�}�Wϸ�&����g��C1�����9�
�b�3��m�(��E�ƭ�l��D�����f�d��f�l�W�W���TӁ��l ��h��*���d�e�4�
�2�<����Y����V��C�U���2�%�3�e�1�n����Aù��l��V�����'�6�o�%�8�8�ǿ�&���R��^	������
�!�e�1�0�N���	����l��F1��*���
�&�
�|�w�}�������F���]���%�6�;�!�;�:���DӇ��P�V ��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�e�3�8�n�}����	����@��X	��*���u�%�&�2�4�8�(���
�ߓ�@��G��U���;�_�u�u�w�}�W�������9��1��*��
�%�6�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���T��Q1�����3�
�m�
�'�>�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�%��(߁�&����lW��h�����!�i�u�'���(���&����V��G1�����4�
�!�'��8�L���YӁ��l ��h��*���d�e�<�
�;�5�(���DӀ��K+��c�����9�<�9�
�c�/���O���F��G1��E���f�3�
�m��3����&��� ��O#��!���!��9�<�;��@�������l�N�����e�3�f�3��e�(�������Z�G1�����<�
�<�n�]�}�W������lV��hZ�� ��b�4�
�0�6�.��������@H�d��Uʲ�%�3�e�3�c�;�(��&����V9��D��*���6�o�%�:�2�.�����ƭ�l��h�����
�!�e�3�:�d�W���&����U9��Q��Mڊ�%�1�;�y�6�����
����g9��_�����e�_�u�u�2�4�}���Y���Z �F��*���&�
�:�<��}�W�������]�F��*���&�
�:�<��}�W���
����@��d:�����3�8�l�u�9�}��������]��[����h�2�%�3�g�;�D���&����R��X ��\���'�}�%�6�9�)���������D�����
��&�d��.�(��P����[��=N��U���u�u�u�'���(���&����Q��G1��U��4�
�:�&��2����B���F����ߊu�u�u�u�w�}����&ù��9��h_�*���6�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=N��U���
�
�
�
��(�F�������R��S�����
�
�
�
�"�l�@���&����G9��h�����0�n�u�u�0�-�����ғ�F9�� 1��*���<�1�f�i�w��(�������]9��PUךU���'�
�
�
�����N����f��T��*���h�3�
�:�2�)����/����`!��D�����'�2�`�d�]�}�W���&����U9��Q��M݊�;��0�6�9��W������W��R��&���7���&�4�4�F�������P��N�����3�e�3�a�1��O؁�����A��C1�I����;�1�
�2�0�$�������l��A��*؊�0�
�d�n�]�}�W������F9��1��U���<�;�%�:�2�.�W��Y����A��B1�@���
�&�<�;�'�2�W�������@N��h��*���$��
�!��.�(������F��h��*���$��
�!��.�(������T9��R��!���d�
�&�
�{�<�(���&����l5��D�����m�u�%�&�0�>����-����9��Z1�\���u�7�2�;�w�}�W��������T�����2�6�d�h�6�����
����g9��1����u�'�;�!��-��������Z��S�����|�u�'�}�'�>��������lW������6�0�
��$�e����N�ƣ�N��h�����:�<�
�u�w�-��������`2��C_�����l�u�'�}�'�>��������lW������6�0�
��$�d����A�ƣ�N��h�����:�<�
�u�w�-��������`2��C_�����d�|�|�!�2�}�W���Y���F��E�� ��`�6�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƫ�C9��h_�*���i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9lǻN��Xʲ�%�3�
�l��m�����Ƽ�\��D@��X���u�2�%�3��d�(�������]9��X��U���6�&�}�
�������ƪ�l��{:��:���g�
�
�0��e�[Ͽ�&����P��h=�����3�8�d�u�'�.��������l��h��*���u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w�-��������`2��C[�����|�u�=�;�]�}�W���Y���T��Q��Lߊ�e�i�u�
���������F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���2�%�3�
�n��G��Y����~3�� ����
�
�0�
�o�f�W���Y����_��=N��U���u�u�u�'��(�F���	���D��o6��-���������/���!����kD��N��U���0�1�<�n�]�}�W���Y����V��=dךU���x�2�%�3��d�(������]F��X�����x�u�u�2�'�;�(��&�ד�@��Y1�����u�'�6�&���(�������F�� 1�����<�y�4�
�>�����*����9��Z1�U���&�2�6�0��	��������l�N�����u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���L����lR����ߊu�u�u�u�w�}��������l��S��*݊�
�;�&�2�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�=�9�W�W���Y���F��G1��*��
�d�i�u���(���
����F�N�����u�u�u�u�w�}�WϹ�	����_��G_��H���������/���!����k>��o6��-���_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������l��V�����'�6�&�{�z�W�W�������lW��h�����2�
�'�6�m�-����
ۇ��P�V�����&�$��
�#�����UӇ��@��T��*���&�`�3�8�c�}��������B9��h��*���
�|�u�u�5�:����Y�����F�����;�!�9�2�4�l�JϿ�&���R��F��*���&�
�:�<��}�W���
����@��d:��݊�&�
�|�:�w�<�(���
����T��N�����<�
�&�$���ځ�
����	�������!�9�2�6�f�`��������V��c1��C���8�`�|�|�#�8�W���Y���F�	��*���d�l�6�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���T��Q��Lӊ�0�i�u�%�4�3��������l�N��Uʰ�1�<�n�_�w�}��������@]ǑN�����3�
�l�
�g�a�W���&����9F�	��*���d�l�%�u�j�-�@�������T]ǻN�����
�
� �g�c�-�W��	����9��Q��Gڊ�d�g�u�u�w�2����I��ƹF��X��*���g�a�%�u�j�-�!���&����lT��h�F���:�;�:�g�~�W�W���&����lW��h��F���%�u�h�_�w�}�W���	����@��A\��Eʢ�0�u�!�%�1��Eف�K���F�G�����_�u�u�u�w�2�(���&���� R��UװU���x�u�
�
��-��������TF��D��U���6�&�{�x�]�}�W���&����l��h�����4�&�2�
�%�>�MϮ�������h/�����1�u�
�
��-����	����9F����ߊu�u�u�u�1�u��������_	��T1�Hʥ�e��4�
�;�t�W������F�N��Uʥ�e��4�
�;��������C9��v1��*���n�u�u�u�w�8����Y���F�N��*ڊ�
�%�#�1�>�����DӖ��l'��G1�����0�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϮ�I����]9��PN�����u�'�6�&�y�p�}���Y����r9��h��*���<�;�%�:�w�}����
�μ�9����*���'�2�u�
���������F��P��U���u�u�<�u��-��������Z��S��*ڊ�
�%�#�1�~�)����Y���F�N��*ڊ�
�;�&�2�k�}�(߁�B���F����ߊu�u�u�u�w�}�(߁�&����Z�
N��E���%�0�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}���&����\�
N��*���0�!�'�
��<����&����Z9��E��@��_�u�u�x�w��B�������R��[
�����;�%�:�0�$�}�Z���YӖ��9��T��*���#�1�4�&�0�����CӖ��P�������2�%�3�e�1�i����AĹ��l��RB�����2�6�0�
��.�Fށ�
����l�N�����u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���H����lW����U���}�4�
�:�$�����&���T��Q1�����3�
�m�
�'�9����P�Ƹ�V�N��U���u�u�%�d��8��������WF������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�%�d��8��������WF������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��Z�����9�
�;�&�0�<����Y����V��C�U���%�d�8�-�6���������l��^	�����u�u�'�6�$�u�(ށ�����l��N��D���-�4�
�9��/��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h_�����%�#�1�|�#�8�W���Y���F���*���
�%�#�1�>�����DӖ��l��h�����_�u�u�u�w�1��ԜY���F�N��D���-�4�
�9��3����E�Ƽ�9��O1��*���
�'�2�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����^��^ �����&�<�;�%�8�8����T�����h��*���&�2�4�&�0�����CӖ��P����*���y�%�d�8�/�-���	�ד�R��G1���ߊu�u�0�<�]�}�W���Y�����T�����2�6�d�h�'�l��������WO�C��U���u�u�u�u�w�-�F�������@��S��*ۊ�4�n�u�u�w�}����Y���F�N��U���
�4�
�;�$�:�K���&¹��K9��R	�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�%�e�����&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��g�����%�#�1�<��4�(�������A	��N�����&�%�g��%�2�(������C9��g�����%�#�1�%�2�t�W�������9F�N��U���}�4�
�:�$�����&���C9��g�����%�#�1�|�#�8�W���Y���F���*���<�1�4�
�;��������C9��g�����%�#�1�_�w�}�W������F�N��U���%�g��'�8���������@��S��*؊�0�<�1�4��1�(������F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C�����'�:�
�9�.�Ͽ�
����C��R��U���u�u�%�g��/��������l��^	�����u�u�'�6�$�u�(݁�����F��1�����
�'�2�u����������E
��=N��U���<�_�u�u�w�}��������]��[����h�%�g��%�2�(��������YNךU���u�u�u�u����������@��S��*؊�0�<�1�_�w�}�W������F�N��U���%�g��'�8��������C9��g�����'�2�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�(ہ�&����]��h^��Hʲ�%�3�e�3�c�;�(��&����V��Y1����u�x�u�
����������l��A�����2�u�'�6�$�s�Z�ԜY�Ƽ�9��c�����
�
�%�#�3�<����&����\��E�����%�6�y�2�'�;�G���M����^��V�����u�%�&�2�4�8�(���
����U��^��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����W��D��E���;�u�:�}�6�����&����P9��
N�����e�3�a�3��e�(�������O�C��U���u�u�u�u�w�-�C���-����T9��1��*���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���&ǹ��g��Y	��*ڊ�%�#�1�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװU���%�a� ��:�3�(���Y����A��h^��*ފ� �d�b�4��8����H��ƹF�N��A����8�;�
������Ӈ��Z��G�����u�x�u�u�'�i�"�������V9��V�����&�<�;�%�8�}�W�������R��RB�����
�
�
�
�"�l�@���&����F��h��*���$��
�!�f�;���P�����^ ךU���u�u�3�}��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�l�(���&���R��Y��]���6�;�!�9�0�>�G������lV��hZ�� ��b�4�
�:�2�t�^Ϫ���ƹF�N��U���
�
�
�<�>�:��������WF������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�%�a��	����&����R��[
��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F���*���%�#�1�<��4�W�������A	��D�X�ߊu�u�
�
��-��������T9��D��*���6�o�%�:�2�.����;����E
����*���%�#�1�%�2�t�W�������9F�N��U���}�4�
�:�$�����&���C9��u1��*���|�u�=�;�]�}�W���Y���C9��u1��*���
�;�&�2�k�}�(ځ�&����_��N��U���0�&�u�u�w�}�W���YӖ��l$��G1�����
�<�u�h�'�h�5���&����C��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�`��4�(���Y����T��E�����x�_�u�u���(���
����@��Y1�����u�'�6�&���(��	�ӓ�l��PB��*ߊ�
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l$��G1�����!�0�u�u�w�}�W���YӖ��l$��Y1����u�
�
�n�w�}�W�������9F�N��U���u�
�
�
�9�.���Y����q9��R	�U���u�u�0�1�>�f�}���Y����C��R�����u�%�c���0����&�����h��*���
� �d�b�6���������9F�C������8�;���(�������@��YN�����&�u�x�u�w�-�A���-����T9��1��*���
�&�<�;�'�2�W�������@N��h��U���
�
�
�
��(�F�������]�V�����&�$��
�#�l����H��ƹF��R	�����u�u�u�3��u��������\��h_��U���6�|�4�1��-��������Z��S�����2�6�0�
��.�Fށ�
����F��SN�����%�6�;�!�;�:���DӁ��l ��h��*���d�b�4�
�8�8�^�������9F�N��U���u�
�
�
�>�4����I����E
��S�����;�!�9�2�4�l�}���Y���V
��d��U���u�u�u�%�a��#�������9��h��U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƹF��hX��*���<�2�0�d�k�}����&ù��9��h_�*���'�!�'�
�l�W�W���TӖ��l0��^�����d�4�
�9�w�.����	����@�CךU���
�
�
�<�>�:��������W9��D��*���6�o�%�:�2�.�����ƫ�C9��1��A���
�m�
�%�3�3�[Ͽ�&����P��h=����
�&�
�e�]�}�W������F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�d�3�8�f�t�������R��X ��*���<�
�u�u�%��(߁�&ǹ��lW��h�����|�|�u�=�9�W�W���Y���F��1��!���;�
�
�
�'�+���Y����\��h�����n�u�u�u�w�8����Y���F�N��*܊�
�<�<�2�2�l���������T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����p9��h��*���&�2�4�&�0�}����
���l�N��B���4�
�9�
�9�.����
����C��T�����&�}�
�
��-����Y����p9��h��*���2�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`����:����E
��N�����u�u�u�u�w�}����:����E
��^ �����h�%�b��6����Y���F��[�����u�u�u�u�w��(���	����l��D��I���
�
�
�%�!�9����B���F���U���u�u�u�0�3�-����
��ƓF�C��*݊�
�;�&�2�6�.��������@H�d��Uʥ�b��<�
�>���������PF��G�����%�b��u���(����Ƽ�9��V�����u�u�7�2�9�}�W���Yӏ��N��h�����:�<�
�u�w��(���	����O��_�����u�u�u�u�w��(�������Z�G1��6�ߊu�u�u�u�;�8�}���Y���F�G1��6���
�<�u�h�'�j�4�����ƹF�N�����3�u�u�u�2�9��������9F���*���<�<�2�0�g�a�W���&����U9��Q��M݊�%�'�!�'��f�}���Y����l^��h�����0�e�4�
�;�}����Ӗ��P��N����u�
�
�
�>�4����I����E
��V�����'�6�o�%�8�8�ǿ�&���T��Q1�����3�
�m�
�'�9�������T9��R��!���d�
�&�
�g�W�W�������F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�d�3�:�l�^Ͽ�ӈ��N��h�����:�<�
�u�w�/�(���&����U��Y�����;�|�|�u�?�3�}���Y���F�G1��"���8�;�
�
��-����E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���
�
�<�<�0�8�G���&����[��G1�����9�2�6�e�]�}�W���Y����Z ��=N��U���u�'�6�&�l�W�W���&˹��G��Y	��*���h�2�%�3�g�;�C���&����R��R�����_�u�u�x�w��(�������l��h�����4�&�2�u�%�>���T���F��1�����;�
�
�
�'�+����
����C��T�����&�}�%�6�{�:����I����l ��V�����:�0�u�%�$�:����&����GW��Q��D���u�u�7�2�9�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��_�����e�u�;�u�8�u��������_	��T1�Hʲ�%�3�e�3�c�;�(��&����\��G�����u�u�u�u�w�}�WϮ�A����Z��P1��D���
�9�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�Ƽ�9��C�����
�
�%�#�3�a�W�������l
��^��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠu�u�%��$�1�(�������9��R��]���4�g�&�3��o�(��J�ƨ�D��]�U���8�
�
�
�"�n�G���P���F��e�����
� �f�e�'�}�J���	����@��A_��E��9�6��3��o�(��B�����V�����
�g�
�d�k�}�(߁�&����Z��N�����g�<�<�<�4�.�(�������P��G]��H�ߊu�u�u�u�'�>��������V��@��U¡�%�<�<�<�e����M����O�I�\ʰ�&�u�u�u�w�}��������_��h_�N���u�'�!�<�>�4����Lù��Z�=N��U���u�%�6�;�#�1�Fځ�I����[����*���
�
�e�3��i�(��I���W����ߊu�u�u�u�'�>��������R��d��Uʦ�9�!�%�
��(�E���	���N��G1�����3�
�f�
�e�%�Ͽ�&����G9��1�N���u�&�9�!�'��(���K�Г�F�F����
�
�
�
�"�o�O���Y����@��C��*��� �g�e�%�~�W�W�������CP��h��F���%�u�h�w�u�*��������f*��Y!��*���<�
�%�,�2�;�(��&�����T�����d�
�a�e�w�1����[���F��[1��݊�
� �f�e�'�}�J���[ӑ��]F��d1�� ���;� �
�e�>���������_��G]��U���6�;�!�9�f��G�������V�=N��U���
�8�m�<�1��Nف�K�����h��C���3�
�m�
�e�2�W���&����l��B1�E���|�_�u�u�2�����&����T��N�U���u�u�u�'�#�4��������9�������8�
�
�
��(�E���	����[�I�����u�u�u�u�w�<�(���
����S��^�U���!�%�d�<�1��A߁�J�����h[�����`�
�f�s�'�m�G߁�&����lU��h�N���u�!�%�f�>�;�(��&���F�N�����&�2�0�}��%�"�������V��Y1�����d�3�
�e��o�W���������T�����d�
��|�2�.�W��B�����hZ�����a�
�f�i�w�}�W���YӇ��P	��C1��M���u�=�;�}�:��(�������l��G��U��|�0�&�u�w�}�W�������]��[��E�ߊu�u�8�
�����I����[�L�����}�<�;�1�1��:���K����lT��^ �����
�
� �f�o�-�^��
����WN��h�����#�m�d�|�2�.�W��B�����h[�����`�
�f�i�w�}�W���YӒ��lR��Q��Aڊ�f�"�0�u�#�-����KŹ��V�
N��R���9�0�_�u�w�}�W���&�Փ�F9��1��N���u�!�%�b��(�D���	��� ��O#��!ػ� �
�e�<��%�(���&����^��F�X��1�"�!�u�~�W�W�������l��h�� ��m�%�u�h�u�� ���Yۊ��l0��B1�A���u�u�%�6�9�)����?����_��^�����u�8�
� �d�k����D�θ�C9��^1��*��
�g�:�u�:��(�������l��d��Uʡ�%�<�<�<�e����M����[�L�����}�:�
�
��(�E���	���R��X ��*���f�e�u�9�2��U�ԜY�Ƹ�C9��^1�����f�
�g�i�w�l�W����Π�P9��Q��Gފ�a�h�4�
�8�.�(���&����_��^�����u�0�4�n�