-- � 2012 National Instruments Corporation.
encrypted
�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�p�}��?����(��G	��4����'�0�&���G������K��B�����0�u�:�2�]�p�8�������c��R��Uʙ�u����0�/�}��=����W��z��G��X�x�X�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T����K�TG��E���%�'�2�#������ƅ�@��Z��ʖ�'�:�4�<�9�W�Zϟ�Ӵ��[��e�����X�x�u�4�>�3�ϗ�
����V��'�����9��3�'�6�4��ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����_�x��'�8�8�z��Y������B�����!�&�=�'�2�.����Y����R��[
�����3�6�u�<�?�3�W���������R�����,��!���}�}��Y����C��Z�����0�u�&�4��1�W���ӄ��Q��[����� �0�!�0�8�8��������\��Y��U���=�;�9�{�]�p�}��>����Z��:d�U����!��1�?�W�Z���Y����G	��[N�����<�!�u�3�6�1����Y����_��U�����0�!�!�{� �}��������VF��[N�����&�!�4�u�'�+�Ϫ�����AF����U���u�0�0�u�9�4�����Ƥ�]��:d�Uʡ�0�u�<�=�#�4�W���	����GH��CаX���:�!�o�_�z�}�4���s���F��V�����:�0�&�4�2�}��������_	����ʔ�u�0�0�4�2�}����W���>l�N��'���!�_�x�u�w���������F��R��[ʆ�;�0�"�u�>�1����
����A	��B�����u�:�u�0�2�<����������@��U���:� �0�&�9�5�����ƾ�@��Q�����0�&�X�x�Z�p�W���<����VF�=C�U���u�;�7�0�$�:��������G	��g'�����u�9�6�u�9�?��������F��C�����0�<�u�0�3�*�����ƅ�z(��DN��ʰ�4�9�1�X�z�P�Z���Y����@��[аX���u�u��1�4�)�W�������Z��DN��ʳ�'�!�!�8�w��9Ϸ�Y����_��:�����0�!�!�0�"�8�����ƭ�l��S�����2�;�'�!�3�?����t���9K�N�����;�_�x�u�w�}�����ƥ�C��Q��U���%�0�u��]�p�W�ԑT����z��C8�����X�x�u�u�w��������� ��ZN�����'��X�x�Z�p�W���+����z��C��U���4�
�:�0�$�:��������V��V��U���6�{��;�2�4�W���	����Z��T��Yʡ�0�0�<�u�8�<�(����ƿ�T�������'�!�1�7�8�6�W�������G	��D�����;�u�<�;�;�W�Z�ԑT����w��x�����u�u�u� �3�8�W���ӕ��GF��	�����0�u�9�6�Z�p�z��Y�Ư�]��a�����X�x�u�u�w�<�(���Y������P�����1�7�:�>�]�p�}��YӅ��R��BаX���u�u��4�.�;�Ϸ�	����\��E������_�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��t����A�����ؠu� �0�<�2�s��������W����N�ߊu�&�u�0�2�3����������c׷���<�,���0��#�������@0��h\�Fʼ�X�u�u�2�9�/��ӶY���F�N�����<�!�u�u�9�8����D����9F�N��U���|�X�u�u�'�/�W���s���F�N�����u�u�u�u�w�}�MϷ�Y����_	��TUаU���u�u�u�u��.����Y���F������9�2�6�X�w�}�W���Y�Ư�]��RN��U���u�u�u�;�$�9������ƹF�N��Uʶ�<�&��9�w�}�W���Y����G��X	��N�ߊu�u�u�u�w�>�������F�N����!�
�:�<��8����Q����R1��C��U���;�:�e�n�]�}�W���Y����z��C8�����u�u�o�<�w�)�(�������F�N��U����4�,�;�w�}�W���Cӏ����h����_�u�u�u�w�}��������F�N��Oʺ�!�u�!�
�8�4�(������X"��V9�����u�:�;�:�g�f�}���Y���F��~ �����<��!�u�m�2��������T��:d��U���u�u�u��6�$����Y���\��B�����9�2�6�n�]�3�W���	����g/��V������g�d�n�]�W��������A��R�����9�:�u�<�'�<�6���1����@��s1�D���&�_�u�u�>�3�Ͻ�����V�N����9�2�6�o�w�l�L�ԜY�ƿ�T������� ��6�o�$�9�������W�:d��Uʦ�2�4�u��'�)����5�����h����_�0�<�X�w�}�%��� ����@��Y�����'�6�&�}�;�t�}���Y����]kǻN��U���3�'�&�;��9�ǝ��Ƹ�V��N��U���u�u�<�u��.����^�Ƹ�V��N��U���u�u�u�u�4�8�������W�:d��U���u�u�u�0�$�;�������A��_�����u�u�u�u�w�}�W�������TF������ ��6�X�w�}�W���Y����]��QUаU���u�u�0�1�>�f�}���Y����C��R��x�ؠu�u�6�4�6�(�W��Y����R/��:d��U�ؠu�u�6�;�"����������G������u�;�u�8�}�1��������������0�n�_�_�w�}�Zϝ�
����\F��CN�����3�'�<�%�#�g�������A��NN��ʼ�%�!�4�u�%�+���������� �����!�4�u�=�$�>����Y����U��CN���ؠu�u�6�0�3�����E�Ư�V��~ �����:�u��%�#�<����Y����P4��S�����'�6�<�&��1�L�Աs���P4��S����u��4�,�"���ӶY���9F������4�<��!�k�}�>�������W*��cךU���_�;�u�0�6�4����t��ƴF��x-��0�������w�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���X�X�x�#�4�3�5���ӧ��#��[��U���6�X�x�#�4�3�Tϟ�Y����XF��X�����<�{�_�x�$�<�W���t����@��+��U���u�-�9�<�w�1��Ӷt���p*��|N��2���u������W��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�ؠX�x�#�6�9�����8����_	��-��x���#�6�;�v��6��������WF��P ���߇x�&�4�u�}�W�Z����Ɖ�WF��S-�����9�X�X�x�w��2���!����r2��y=��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T����>l�A��ʗ�2�;��1��-����+����>l�A�����&�4�1�'�w�4����Y����[��X�����!�_�x�&�6�}�%������E��YN���ߧ_�x�����0���Y����p'��x ��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�Ӷt����@��,�����1�u�-�9�>�}�������E��YN�����'���<�w�1�W������9K��D��U���_�x�&�4�w�3�W���Y����R��x�� �ؠX�x�u���	�8���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s��