-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǶd�����,�<�0�n�]�.�W���ݕ��l
��^��D��4�9�u� �2�4��������T��B �����{�9�n�_�9�4�ϳ�I����uV��1�����d�a�
�4�w�.�}���Y����A��=N��U���u�u�u�0��$����Y�ƿ�A��T��W���6�w�u�u�w�}�W���Yӂ��W��N��Oʼ�!�2�'�o�w�o�W���Y���F������u�u�o�<�#�:���Y���F�N��U���8�8�&�/�w�}�MϷ�����\�d��U���u�u�u�%�%�}�}���Y���F��S�U���o�<�u�!��2����������S��Dʱ�"�!�u�|�w�}�W���Y����VV�N��U���;�&�1�9�0�>�W���Y���F��N��U���u�u� �u�#�����&����\��@����1�"�!�u�~�W�W���Y���R��N��U��<�u�!�
�8�4�(�������D��_C����!�u�|�u�w�}�W���YӅ��F�N��U���&�1�9�2�4�}�W���Y�����N��U���u�;�&�1�;�:��������W��C��U���;�:�e�n�]�}�W���Y�ƻ�F�N��Oʼ�u�!�
�:�>�f�}���Y���F��\N��U���u�u�;�&�3�1����s���]�R �����!�n�_�_�%�5��������G
��QN��E��`�e�
�
�"��(��@������=d�����u�1�'�
�:�}�W���&����P9��T��]���1�=�d�1� �)�W���Y����VF��Z1�����<�u�'�4�w�m��������I�N��U���
�:�<�
�2�)��������W��X����n�_�=�'�3�+�����ƾ�^F��Z�����,�_�4�!�>�(�ϭ�����@��RN����;�n�_�!�%�?���� ����^��[��ʧ�8�o�#�'�6�1�W���[����X9��ZL����<� �0�'�:�.����Cӕ��Z��=�����!�u�4�
�#�1�W��������^��ʼ�u�0�
�,�2�W��������v7��a/��;���������!���Cӕ��Z��=d�����_�_�0�:�.�<����&����W9�������u�4�1�e�w�?����Y�����E^�����h�4�1�e�]�p��������G��D�����3�u�u�u�>�}�4���&����t#��V
��E���u�0�
�<�2�l�W������F�N�����e�!�%�i�w�2����Y���A�=N��U���9�0�_�u�w�}�W�������l��R�����e�_�u�u�w�3�W���s�˿�]��D�����&�4�0�:�]�3�W�������9l��Z�����6�0�&�e�w�/����Yۅ��F�U���ߊu�u�3�}�;�z����Y����P
��
N��R���=�;�u�u�w�}�������A��N�����u�u�u�u�w�}����DӔ��%��a1��!����4�1�e�#�-�^���Y���F��Y
���ߊu�u�;�u�1�W��������@]Ǒ=�����,�4�6�&��g�������P
��N�����u�u�u�<�w�>�Ȼ�����]��[��U��|�!�0�_�w�}�W����ί�F�_��U���;�_�u�u�w�}�W����λ�F�_��U���;�_�u�u�w�}�W���Y�ƾ�^N��y8��;����}�1�'�~�}�JϺ�B���F�N��Uʰ�1�<�n�u�w�}�Wϻ�ӏ��9F���U���_�;�u�'�4�.�L�Զ����G
��=d�����,���n�"�8�>���W����_	��T1�C���9�n�_�;�>�$���N�ӊ�U9��U��E��a�u�&�u�w�:������ƹF�N�����<�!�u�u���2���D����9F�N��U���'�&��;�2�g�>���>���F��=N��U���u�1�'�&� �9���0����v4�
N�N���u�%�'�u�]�}�W���Y����GF��~ ��!�����n�u�w�}�WϽ�����}F��s1��2���_�u�u�u�w�9����I����}F��s1��2������}�3�/�������W��x9��:��n�u�u�u�w�>�G��0�Ɵ�w9��p'�����u�u�u�e�m��#ύ�=����z%��r-��'�!��1�=�z�l�3���-����l�N��Uʴ�1�0�&�u�w��$���5����l0��c!��4���0�&�<�!�w�}�W���7���]ǻN��U���0�u�u����;���:���F�N��D���u��
���L���Y�����N��U���
���
��	�%ǚ�����G�_��:����e�|�_�9�}���� ����A��C�� ���4�6�u�3�:�m�@���I����Q��1�A���&�u�u�6�:�2��������S��Q1�����e�d�a�
�6�}����Y�����CN��U���u�u�u�u�4�6�Mϗ�Y����)��tUךU���u�u�u�u�3�/�W���7ӵ��l*��~-��0����_�u�u�w�}�W�������z(��c*��:���n�u�u�u�w�}�Wϯ�Y�ƃ�gF��s1��2������n�w�}�W���Y����W��T��;ʆ�������8��Y���F�N�����u������4�ԜY���F�N��U���������!���6��ƹF�N��U���0�u�u����;���:��ƹF��Y
�����;�;�n�_�]�8��ԜY�ơ�_��(��*ڊ� �
�
�g�n�/����C�Ư�^��R ����b�`�e�
��(�(߁�K�ߓ�RǻN�����8�%�}�u�w�}�WϽ����P
��=N��U���u�1�'�u�i�<����
��ƹF�N�����k�6�e�_�w�}�W���I���BV�N��U���4�1�d�h�w�9����H���F�N��D��u�0�y�u�w�}�WϺ�Y����JǻN��U���0�u�k�"�f�f�}���Y����Z��C��N�ߠ