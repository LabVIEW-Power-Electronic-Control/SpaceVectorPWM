-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�������(���
����GF�N�����9�u�u����;���:���F��h��U���������}���Y����G��T��;ʆ�����]�}�W�������	F��cN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�%�<���6����g"��x)��N���u�<�
�9�?��(���Y����g"��x)��*�����}�d�3�*����P���F��h��*؊�u�u�����0���/����aF�N�����u�|�_�u�w�3����&ù��	F��=��*����
����u�FϺ�����O��N�����0� �;�e�m��#ύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����V��Y1�Oʚ�������!���6���F��@ ��U���_�u�u�%�%�)����Y�ƃ�gF��s1��2������u�d�}�������9F������'�
�u�u��}�#���6����e#��x<��Bʱ�"�!�u�|�]�}�W�������z(��c*��:���u�n�0�1�]�W��������A��R��U���8������(���Y���F�T�����u�%�6�;�#�1����H����g"��x)��U��r�r�_�u�w�2����Ӈ��P	��C1�����e�o�����4��Y���9F������!�4�
��$�l����I����g"��x)��*�����}�u�8�3���Y���V��L�U���6�;�!�;�w�-�$�������^9��N��1��������}�CϺ�����O�
N��E��w�_�u�u�8�.��������l��h��*���u��
����2���+����W	��C��\��u�e�d�e�l�}�WϽ�����GF��h=�����3�8�f�o���;���:����g)��Z�����:�e�u�h�u�l�G���s���P	��C��U����
�!�
�$��W���-����t/��a+��:���a�1�"�!�w�t�M���H����]ǻN�����4�!�4�
�8�.�(���K���5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��2����¹��	F��s1��2������u�g�9� ���Y���F�UךU���:�&�4�!�6�����&����lW�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��_�����u�:�&�4�#�<�(���
���� T��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�:�&�6�)��������_��h]��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�D���_�u�u�:�$�<�Ͽ�&����G9��Y��L��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�e�d�g�l�F��H����F�T�����u�%�6�;�#�1�D݁�<����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��I����]ǻN�����4�!�4�
�8�.�(���K���5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����W�=N��U���&�4�!�4��2�����ԓ�\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����W��UךU���:�&�4�!�6�����&����lV�=��*����
����u�DϺ�����O�
N��E��e�e�e�e�g�f�W�������R��V�����
�#�g�d�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��I����V��^�E��e�e�e�e�f�l�U�ԜY�Ư�]��Y�����;�!�9�f���1���?����g"��x)��*�����}�d�3�*����P���V��_�D��d�d�d�d�f�l�F��H����]ǻN�����4�!�4�
�8�.�(���K����V��N�&���������W��Y����G	�N�U��e�e�e�e�g�m�G��I����V��^�E��u�u�6�;�#�3�W�������l
��1�Oʆ�������8���J�ƨ�D��^��O���e�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[�*��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D������o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�d�d�n�w�}��������R��X ��*���g�d�u�u���8���&����|4�_�����:�e�u�h�u�m�G��I����V��^�E��e�e�d�e�u�W�W�������]��G1�����9�f�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�E��e�e�e�d�g��}���Y����G�������!�9�d�
�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��UךU���:�&�4�!�6�����&����lW��N��1��������}�D�������V�S��E��e�e�e�e�g�m�G��I����V��^�N���u�6�;�!�9�}��������EU��+��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��_�D���_�u�u�:�$�<�Ͽ�&����G9��1�Oʆ�������8���Kӂ��]��G��H���d�w�_�u�w�2����Ӈ��P	��C1��A���o������!���6�����Y��E���h�w�d�d�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�g�m�U�ԜY�Ư�]��Y�����;�!�9�g�g�g�$���5����l0��c!��]���:�;�:�e�w�`�U��B�����D��ʴ�
�:�&�
�!��W���-����t/��a+��:���g�1�"�!�w�t�M���H���9F������!�4�
�:�$��܁�Y�Ɵ�w9��p'��#����u�g�1� �)�W���C���V�=N��U���&�4�!�4��2�����Г�u ��N��1��������}�F�������V�S��E��d�d�d�d�f�l�U�ԜY�Ư�]��Y�����;�!�9�d��m�G��*����|!��h8��!���}�`�1�"�#�}�^��Y����V��^�E��e�n�u�u�4�3����Y����\��h��F��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I��ƹF��X �����4�
�:�&��+�(���Y����)��t1��6���u�g�1�"�#�}�^��Y����]ǻN�����4�!�4�
�8�.�(���&����`2��{!��6�����u�g�3�*����P���V��UךU���:�&�4�!�6�����&����F��d:��9�������w�o��������\�^�W�ߊu�u�:�&�6�)��������_��N�&���������W������\F��T��W��w�_�u�u�8�.��������]��[�*��o������!���6���F��@ ��U���o�u�e�e�g�m�G��I����V��^�E��e�e�n�u�w�>�����ƭ�l��D��ي�u�u��
���(���-���F��@ ��U���o�u�e�e�l�}�WϽ�����GF��h�����#�d�f����W���-����t/��a+��:���f�u�:�;�8�m�W��[����W��_�D��d�d�d�d�f�l�F��B�����D��ʴ�
�:�&�
�!�l�C��I����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��2�����ԓ�F��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-��������lU�=��*����
����u�W������F��L�W�ߊu�u�:�&�6�)��������_��hZ��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�:�$�<�Ͽ�&����G9��1�Oʆ�������8���Jӂ��]��G��H���e�d�n�u�w�>�����ƭ�l��D�����e�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�e�w�_�w�}��������C9��Y����
�e�e�e�g�g�$���5����l0��c!��]��1�"�!�u�~�g�W��H����V��^�E��e�e�e�e�g�m�U�ԶY����Z��[N��*���3�8�o����0���/����aF�
�����e�u�h�w�g�m�U�ԜY�ƭ�G��B�����0�6�1�;�w�}�������F��C�� ���3�8�0�6�3�3�W�������l ��T�����9�<�u�;�9��}���Y����R
��G1�����0�
��&�f�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������	F��x"��;�ߊu�u�<�;�;�.��������lW��N�&���������W������\F��d��Uʦ�2�4�u�
�6�o�E���&����CT�=��*����
����u�FϺ�����O��N�����4�u�
�4�e�o����H����	F��s1��2������u�d�}�������9F������;�"�<�;�>����H����	F��s1��2������u�g�9� ���Y����F�D�����0�&�2�7�#�/���H����`2��{!��6�����u�e�3�*����P���F��P ��U���
�
� �g�n�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��*���
�m�b�o���;���:����g)��^�����:�e�n�u�w�.����Y����Z��D��&���!�
�&�
�w�}�#���6����9F������4�
�<�
�3��O��;����r(��N�����4�u�8�
��8�(��A����g"��x)��*�����}�u�8�3���B�����Y��������!�f�d�!�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�-������&����e9��E��D��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���&�ғ�V��Z�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�;����I����	F��s1��2������u�g�9� ���Y����F�D�����9�
�0�
�o�h�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�����0�8�a�`��;�(��&���5��h"��<������}�e�9� ���Y����F�D�����-�
�:�0�#�/�(��&����T9��^��U���
���
��	�%���Kӂ��]��G�U���&�2�4�u�/��2�������9��Q��Eڊ�g�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�	����K)��h_�*���0�
�m�m�m��3���>����v%��eN��Gʱ�"�!�u�|�]�}�W�������Z��^��*���
�m�m�o���;���:����g)��^�����:�e�n�u�w�.����Y���� _��R	��M��o������!���6�����Y��E��u�u�&�2�6�}�(���K����U�� Z��G��������4���Y����W	��C��\�ߊu�u�<�;�;�-�!���&�Փ�V��Y�Oʆ�������8���H�ƨ�D��^����u�<�;�9�9�*��������U��^��F��������4���Y����\��XN�N���u�&�2�4�w�8��������l��h_�@��������4���Y����\��XN�N���u�&�2�4�w�0�(�������9��T��!�����
����_�������V�=N��U���;�9�!�%�f�����A���5��h"��<������}�w�2����I��ƹF��^	��ʇ�;�0�
�9��3����&����CT�=��*����
����u�W������]ǻN�����9��;�0��1�(���
����lW��N�&���������W������\F��d��Uʦ�2�4�u�4�0�l��������l ��]�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�����&����I��D1����e�u�u����>���<����N��S�����|�_�u�u�>�3�Ϯ�M¹��U��X��G��������4���Y����\��XN�N���u�&�2�4�w��F�������
V��N��1��������}�GϺ�����O��N�����4�u�8�
��(�A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�
�0�
�n�n�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��h��*���$��
�!��.�(���Y����)��tUךU���<�;�9�4��4�(���&���$��{+��N���u�&�2�4�w�(�(������� 9��^�����2�
� �d�g��D��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��X��&���:�
�f�"�>�8��������T9��^��U���
���
��	�%���Y����G	�UךU���<�;�9�'��;�(��N����	F��s1��2������u�d�}�������9F������'��'�2�f�o�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��E1��G���
�e�d�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����A9��1����f�u�u����>���<����N��
�����e�n�u�u�$�:����&����lT��Q��E���%�u�u����>���<����N��
�����e�n�u�u�$�:����&����lT��E��D��u�u��
���(���-��� U��X����n�u�u�&�0�<�W�������lT��Q��E���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϱ�&����9��h��*��d�o�����4���:����V��X����n�u�u�&�0�<�W���&����l ��^�*��o������!���6�����Y��E��u�u�&�2�6�}�����ޓ�V��Z�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)��������
S��N��1��������}�GϺ�����O��N�����4�u�0�
�:�l�(���H����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'�n����H����	F��s1��2������u�g�9� ���Y����F�D�����8�
�f�3��o�@���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����g�
�0�
�n�d�Mύ�=����z%��r-��'���e�1�"�!�w�t�}���Y����R
��G1�����0�
��&�c�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}��������V9��E�� ���`�
�
�
�"�l�Oف�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�!��&��)��������l0��h��*��a�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�/����@9��h_�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������U��[��G��������4���Y����W	��C��\�ߊu�u�<�;�;�)���&����W��N�&���������W��Y����G	�UךU���<�;�9�!�'�n�(���H�ד� F��d:��9�������w�m��������l�N�����u�
� �d�b�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h��*���d�l�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӗ��G9��h_�*��o������!���6�����Y��E��u�u�&�2�6�}����
����9��h\�*��o������!���6�����Y��E��u�u�&�2�6�}�(���K�ד�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�0�(ށ�����l��N��1��������}�D�������V�=N��U���;�9�!�%�1��C܁�K����g"��x)��*�����}�u�8�3���B�����Y��������!�f�j�!���&����CT�=��*����
����u�FϺ�����O��N�����4�u�4�'��(�E���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�
� �g�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h ��*��� �g�f�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������A��P��*���g�m�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӂ��V��h�����
�b�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ʈ�^��RZ�����'�4�
�
�"�o�N���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����'�
� �g�n�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��E����
�
� �f�c�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Y
�����
� �f�e�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W�������	��E�����
�l�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƣ�T9��T1�����
�g�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�CW��B1�M���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������l��B1�C���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'��݁�@����l ��Z�����u��
����2���+������Y��E��u�u�&�2�6�}�(���K����9��h]�*��o������!���6���F��@ ��U���_�u�u�<�9�1����A���� Q��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�3�'��$�������l0��B1�C���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���/����W9��D��*���g�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�C9��d����l��d�3��e�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����m�3�
�f��l�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��Z��E���
�`�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƾ�9��hZ�*��o������!���6�����Y��E��u�u�&�2�6�}�(���K����S��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�$�>��(���M�ғ� F��d:��9�������w�m��������l�N�����u�7�4�&�0��(���M�ғ�F��d:��9�������w�m��������l�N�����u�
�4�g�f����M����	F��s1��2������u�f�}�������9F������!�%�&�3��j�(��Cӵ��l*��~-��0����}�`�1� �)�W���s���@��V��*��� �!�l�3��m�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��'���9�
�
� �b�e����Y����)��t1��6���u�f�1�"�#�}�^�ԜY�ƿ�T����*���3�
�l�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����a��R\�����;�&�3�
�f��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��D؊� �`�e�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������\	��O)��:���d�a�3�
�a��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��U��*���e� �
�c��(�B���	����`2��{!��6�����u�e�3�*����P���F��P ��U���9�-���#�l�O���&����CT�=��*����
����u�W������]ǻN�����9�!�%�f��(�B���	����`2��{!��6�����u�d�3�*����P���F��P ��U���
�:�0�!�%��Oہ�&����
W��N�&���������W��Y����G	�UךU���<�;�9�!�'�i����OĹ��\��c*��:���
�����}�������9F������6�'�,�d�1��Eہ�K����g"��x)��*�����}�u�8�3���B�����Y�����!�1�/�'�$�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʥ�;�!�<�
�"�k�B���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����2�
�d�3��h�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
� �c�c�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������R��*���&�d�3�
�d��D��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��G1�*��� �c�e�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������A��P�*���:�2�;�<��(�A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���d�f�1�8�%�<�(���O�ԓ�F��d:��9�������w�m��������l�N�����u�8�g�3��j�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����9�"�d�3��e�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����:�
�
� �a�l����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����F���
�l�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ʈ�^��R1��ۊ� �c�l�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������]��Q��*ۊ�:�
� �b�f�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h8��G��a�8�-�3��m�(��Cӵ��l*��~-��0����}�`�1� �)�W���s���@��V��*���g�d�d�
�"�j�C���Y�Ɵ�w9��p'��#����u�d�u�8�3���B�����Y�����d�
� �b�f�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��Q�����
�0�8�a�o�����Kʹ��\��c*��:���
�����e��������l�N�����u�6�%�3��e�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����
�e�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G_�� ��d�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������]	��Q��@ӊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&ƹ��lP��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2���������9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�(�������l �� [�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	�Փ�V��P�����b�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����9��hX�*��o������!���6�����Y��E��u�u�&�2�6�}��������lQ��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����&����A��h��B���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϭ�����9��hV�*��o������!���6�����Y��E��u�u�&�2�6�}�����ӓ�F9�� 1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����&����_��N�&���������W������\F��d��Uʦ�2�4�u�0��0�@���&����CT�=��*����
����u�W������]ǻN�����9�&�9�!�'����N����	F��s1��2������u�g�9� ���Y����F�D�����'�6�;�
�"�e�N���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����9�3�
�d��n�Mύ�=����z%��r-��'���g�1�"�!�w�t�}���Y����R
��R��ۊ� �m�`�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����\��X ��*���m�d�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӊ��P	��1��*���
�g�o����0���/����aF�
�����e�n�u�u�$�:�������� 9��hV�*��o������!���6���F��@ ��U���_�u�u�<�9�1�����ԓ�F9�� 1��U����
�����#���Q����\��XN�N���u�&�2�4�w�%�(�������U��a1��*��
�g�o����0���/����aF�N�����u�|�_�u�w�4��������_S��B1�@���u�u��
���(���-��� T��X����n�u�u�&�0�<�W���*����U�� \��F��������4���Y����W	��C��\�ߊu�u�<�;�;�3� ���A����^��G]��U���
���
��	�%���Kӂ��]��G�U���&�2�4�u�2��؁�����l��N��1��������}�D�������V�=N��U���;�9�3�%�9�9�(�������l0��V�����f�
�d�o���;���:����g)��]����!�u�|�_�w�}����ӈ��`��h��L���%�u�u����>���<����N��
�����e�n�u�u�$�:��������
9��hW�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������l��C1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������_W��Q��GҊ�f�o�����4���:����U��S�����|�_�u�u�>�3�ϰ�����W��V�����f�
�d�o���;���:����g)��]����!�u�|�_�w�}����ӈ��`��1��*��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������_W��Q��@ي�f�o�����4���:����U��S�����|�_�u�u�>�3�ϰ�����9��hW�*��o������!���6���F��@ ��U���_�u�u�<�9�1��������l��C1����� �l�l�%�w�}�#���6����e#��x<��Gʱ�"�!�u�|�]�}�W�������V��[_�����b�
�f�o���;���:����g)��\�����:�e�n�u�w�.����Y����V
��h��L���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϰ�����9��hW�*��o������!���6�����Y��E��u�u�&�2�6�}�(���K�ӓ�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w�����M����
T��G]��U���
���
��	�%���Kӂ��]��G�U���&�2�4�u�:��B���&����l��N��1��������}�D�������V�=N��U���;�9�!�%�f����H����\��c*��:���
�����n��������l�N�����u�
�4�g�d�;�(��&���5��h"��<������}�e�9� ���Y����F�D�����
�4�g�g��(�O���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʡ�%�d�
� �f�o�(��Cӵ��l*��~-��0����}�f�1� �)�W���s���@��V�����m�3�
�e�`�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��C��Dӊ� �d�f�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������h[�����e�b�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӏ��CW��B1�@ߊ�g�o�����4���:����V��X����n�u�u�&�0�<�W���	�ӓ�\��B1�Bي�g�o�����4���:����V��X����n�u�u�&�0�<�W���&�ѓ�F9��Y��G��������4���Y����\��XN�N���u�&�2�4�w�8�(���@����V��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2����N����\��Y1��*��d�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CW��h
�����;�3�
�d�n�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����
� �d�d��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���d�g�
�d�m��3���>����v%��eN��Aʱ�"�!�u�|�]�}�W�������^��1��*��e�%�u�u���8���&����|4�Z�����:�e�n�u�w�.����Y����_T��1��*��f�%�u�u���8���&����|4�Z�����:�e�n�u�w�.����Y����@��h]�� ��`�
�a�o���;���:����g)��\�����:�e�n�u�w�.����Y����Z��^��*���d�a�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƽ�]	��^\�� ��c�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����T9��h_�L���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������9��h_�D���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����K����lW�� 1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'�3��������W��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�2�.�����֓�\��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������VU��^1��*��d�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������U
��h\�� ��e�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����U
��h\�� ��m�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����A ��@1�����3�
�g�l�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������R��*���g�3�
�g�d�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��@���
�g�d�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����Q��E	��*���d�g�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������9��h_�L���u�u��
���(���-��� V��X����n�u�u�&�0�<�W���&�Փ�R��Q��G���%�u�u����>���<����N��
�����e�n�u�u�$�:����&����lU��Q��G���%�u�u����>���<����N��
�����e�n�u�u�$�:��������l ��\�*��o������!���6�����Y��E��u�u�&�2�6�}��������lU��B1�M܊�f�o�����4���:����V��X����n�u�u�&�0�<�W�������l ��]�*��o������!���6�����Y��E��u�u�&�2�6�}����&¹��lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�5�0��������lW��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Eہ�����9��T��!�����
����_�������V�=N��U���;�9�%�;�#�e�ށ�����9��T��!�����
����_�������V�=N��U���;�9�;�"�>�3����&����ZW��B1�GҊ�g�o�����4���:����V��X����n�u�u�&�0�<�W�������
9��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������_	��1��*��c�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������_	��1��*��g�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������U
��h]����� �d�`�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����Q��E	�����
� �d�`��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��a��*���3�
�g�g�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��Z��ߊ� �d�c�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����C9��[\��Dي� �
� �d�`��D��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T�������f�g�
� �f�j�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����2�6�0�
��.�B������5��h"��<��u�u�&�2�6�}��������lQ��T��:����n�u�u�$�:��������l��C1��*��e�%�u�u���8���&����|4�]�����:�e�n�u�w�.����Y����_T��1��*��f�%�u�u���8���&����|4�]�����:�e�n�u�w�.����Y����S��B1�GҊ�a�o�����4���:����W��X����n�u�u�&�0�<�W���
����Z��h��D��
�f�o����0���/����aF�
�����e�n�u�u�$�:����&����ZR��B1�FҊ�g�o�����4���:����V��X����n�u�u�&�0�<�W�������U��^�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�?��������U��Z�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����S��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�%�9�)�O���&����P��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�;� �4����&ù��G9��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������VU��^\�� ��b�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����A ��@1�����a�e�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӊ��A ��@1�����a�c�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӓ��V��X��*���
� �d�l��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��Z�����<�
� �d�o��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��G1��؊�g�3�
�a�a�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��U�����
� �d�l��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��a��*��
� �
� �f�m�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��*���g�a�g�
�"�l�F݁�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�!��&��)��������l0��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������G9��D�����!�'�
�g��j����J�ѓ�F��d:��9�������w�n�W������]ǻN�����9�3�%�-��$��������P��X��*��� �d�g�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W������� ��h��6���
�!� �!�%��N�������Q��N�&���������W��Y����G	�UךU���<�;�9�3�'�>�(�������F��E��L���f�3�
�`�c�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��Q�����4�0��'�4�(���&����U��X�����u��
����2���+������Y��E��u�u�&�2�6�}��������V9��E�� ���a�
�
�
�"�l�A؁�J����g"��x)��*�����}�d�3�*����P���F��P ��U���4�g�g�e�1�-���� ����`��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������G9��D�����!�'�
�g��;�(��N����	F��s1��2������u�d�}�������9F������3�%�6�
�6�8�$�������lR��a1�����`�a�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�C9��h-�����'�6� �0�c��(݁�����9��T��!�����
����_������\F��d��Uʦ�2�4�u�-��)�4���&����P��R1�*���
� �d�l��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��h8��G��l��9�
��(�F��&���5��h"��<������}�f�9� ���Y����F�D�����-�
�!��$���������P��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������G9��D�����!�'�
�c��o����O�ғ� F��d:��9�������w�n�W������]ǻN�����9�3�%�6��<��������A��1��F���
�c�d�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����U��T������'�6� �2�h�(���&����T��G]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�:��O���&����l��N��1��������}�DϺ�����O��N�����4�u�8�
�n�;�(��L����	F��s1��2������u�g�9� ���Y����F�D�����8�
�`�3��h�D���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�����g�3�
�c�n�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��h^�F���e�c�
�
�"�l�A܁�J����g"��x)��*�����}�e�3�*����P���F��P ��U���8�<�!�� �4����
����U��Y�����u��
����2���+������Y��E��u�u�&�2�6�}����I����P��h�Oʆ�������8���Jӂ��]��G�U���&�2�4�u�:��F���&����l��N��1��������}�GϺ�����O��N�����4�u�8�
�a�;�(��M����	F��s1��2������u�d�}�������9F������<�8�f�3��k�D���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V��*��f�e�e�b�����IĹ��\��c*��:���
�����m��������l�N�����u�&�8�<�#�� �������Z��1��*��`�%�u�u���8���&����|4�^�����:�e�n�u�w�.����Y����T��B1�G݊�a�o�����4���:����U��X����n�u�u�&�0�<�W���&�Փ�F9��]��F��������4���Y����\��XN�N���u�&�2�4�w�0�(������� S��N�&���������W��Y����G	�UךU���<�;�9�<�:�i����N�ѓ�F��d:��9�������w�m��������l�N�����u�
�g�f�g�m�Oف�&����S��G]��U���
���
��	�%���Iӂ��]��G�U���&�2�4�u�$�0����/����G��D�����3�
�b�l�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��S�����
�'�!�
�$�4����
����lW�� 1��U����
�����#���Q����\��XN�N���u�&�2�4�w�.��������A��h�����g�6�&�
�"�l�E܁�H����g"��x)��*�����}�d�3�*����P���F��P ��U���8�<�!�� �4����
���� 9��D�� ��b�
�d�o���;���:����g)��]����!�u�|�_�w�}����ӈ��`��W�����3�
�f�a�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������y=�����u��
����2���+����W	��C��\�ߠ_�0�<�_�]�W�W���TӒ����E��U���!�u�4�
��;����Ӓ����C�����;�{�x�_�w�}����&����R��P �����o�%�:�0�$�<�(���P�����^ ךU���u�u�3�}�'�>�Ȼ�����]��G1����u�d�|�!�2�W�W���Y���F��F��*���u�u�d�|�#�8�}���Y���F�N������3�8�i�w�-�$���¹��^9��=N��U���u�u�u�9�2�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C��U���u�u�u�u�w�}�W���YӇ��p5��D��Hʴ�
��3�8�]�}�W���Y���F�R ����_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9l�N�U���<�;�%�:�2�.�W��Y����A	��D�����9�|�u�u�5�:����Y����������0�0�!�4�3�<�(���Y���O��_��U���u�u�u�u�>�}�_ǿ�&����G9��P��D��4�
�0�u�9�}��������_	��T1�Hʴ�
�<�
�&�&��(���&����O������u�u�u�u�w�}�Wό�����R
��X ��*���
�m�c�i�w�<��������]��Q��GҊ�g�_�u�u�w�}�W���Y�ƞ�]��h��*���:�
�0�
�n�n�K�������l��h����� �`�a�%�l�}�W���Y���F���*���-� �
�c���(���&����Z�Q��4����!�d�l��n����Lǹ��l�N��U���u�u�u�3�'��0�������l0��R	��M��i�u�-�
��%����Jƹ��U��^��G�ߊu�u�u�u�w�}�W�������W��R��A����'�2�d�b�}�Jϸ�	����V9��E��Eߊ�
� �f�c�'�f�W���Y���F�N�����2�7�!�d�%�:�F��Y����l0��1�*���a�a�%�}�b�9� ���Y���9F�N��U���u�u�u�
�f�4����H����[��hZ�����
�a�
�g�]�}�W���Y���F�G1��؊�f�'�2�d�`�}�JϮ�/����U��B1�A���n�u�u�u�w�}�W���Yӕ��]��h_�����m�m�i�u�/��2�������9��Q��Eڊ�g�f�u�:�9�2�D���s���F�N��U���!�%�d�
�2��O��E�Ƹ�C9��h��A���%�n�u�u�w�}�W���Y����^��1����a�u�h�3�'��$�������l0��h��F���%�}�d�1� �)�W��B���F�N��U���u�8�
�l�%�:�F��Y����K��r)�� ���f�
�
� �c�m����Aӂ��]��V����u�u�u�u�w�}�W���&ʹ��T9��V��Hʼ�
�9�=�
��u�FϺ����� W�=N��U���u�u�u�u�w�1�(���&����Z�B�����l�
�g�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dךU���x�4�&�2�w�/����W���F�G�����}�%�6�>�]�}�W������F�N��U´�
�9�r�#�9�}����	����[�I�����_�u�u�u�w�}�W���Q�έ�l��D�����
�u�u�%�4�t����Q����\��h�����u�u�%�&�0�>����-����l ��h]��\ʡ�0�_�u�u�w�}�W���Y�ƪ�C9��h-�����'�6� �0�b��(؁�����R�
N�����
�4�0��%�>����LŹ��9��h_�C���n�u�u�u�w�}�W���YӒ��lT��E��D��u�h�!�%�e����LĹ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�4�
�:�$�����&���R��^	������
�!�
�$��^Ͽ��έ�l��D�����
�u�u�%�4�t�������R��C��U���%�6�;�!�;�:���P����[��N��U���u�u�u�u�9�*��������T9��^��Hʥ��9�
�
�"�o�B���Q����\��XN�\�ߊu�u�u�u�w�}�W���&����lT��R	��M��i�u�
�4�e�o����Hƹ��l�N��U���u�u�u�&�0�?��������F������&�3�
�a��o�C�������R��d��U���u�u�u�u�w�)��������W��S�����
� �g�l�'�f�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠu�u�x�u�$�4�Ϯ�����F�=N��U���6�&�u�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��R��u�=�;�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1����|�u�=�;�w�}�W���Y���F��E1�����g�
�0�
�n�l�K�������WW��1��*��d�%�n�u�w�}�W���Y���	��h=�����d�
�'�!��.��������
T��S�� ���0�!�'�d��/����
����l ��^�*��_�u�u�u�w�}�W���Y����_T��1����f�u�h�%��1�(�������W��UךU���u�u�u�u�w�}�(���&����_��R�����g�3�
�e�f�-�L���Y���F�N��U���
�0�
�l�b�a�W���&����W��G\�U���u�u�u�u�w�}��������l��h_�@��u�0�
�8�f����I����l�N��U���u�u�u�&�;�)��������
P��S�����8�d�
� �f�o�(��s���F�N��U���&�9�!�%��8�(��A���@��C��*���d�m�
�g�]�}�W���Y���F�C��B���2�d�d�u�j�)��������9��d��U���u�u�u�0�3�4�L���Y����������u�;�u�'�4�.�L�ԜY����� ��ʦ�4�0�}�%�������Ƹ�VF��V�����<�0�u�x�w�}����*����l��^	�����u�u�'�6�$�}����������t=�����4�
�0�_�w�}����s���F�T��U����
�&�u�$�}�W���Y�����YN��*���&�d�3�8�g�`�W���Y���F�N��U���}�}�%�6�9�)���������T�����;�!�}�%�$�<�������]��[����|�|�!�0�]�}�W���Y���F�N������3�8�i�w�-�$�������^9��=N��U���u�u�u�u�w�1����Y���F�N��U���u�%��
�$�}�JϿ�&����GW��D��N���u�u�u�u�w�}�Wϻ�ӏ��9F�N��U���u�=�;�4��	��������[�=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���4�
��3�:�a�W���*���� 9��Z1����u�u�u�u�w�}�W������F�N��U���u�u�u�%������DӇ��`2��C\�����n�u�u�u�w�}�W���YӃ����=N��U���u�u�u�=�9�<�(���
�Փ�@��S����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�4�
��;���Y����g9��1����_�u�u�u�w�}�W���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:��ي�&�
�n�u�w�}�W���Y����������u�u�u�u�w�5�Ͽ�&����GR��D��U��_�u�u�u�w�}�W���Y�����T�����2�6�d�h�6���������F�N��U���u�u�u�u�6��$������R��c1��@���8�a�_�u�w�}�W���Y���V
��=N��U���u�u�u�u�w�}�W���7����^F���&���!�
�&�
�l�}�W���Y���F���U���_�u�u�u�w�}�W���Ӈ��`2��C[�����u�k�_�u�w�}�W���Y���Z ������!�9�2�6�f�`��������[��N��U���u�u�u�u�w�}����*����Z�V��!���d�3�8�e�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y����	��R��H���_�u�u�u�w�}�W���Y����`9��ZN�Uȍ���n�u�w�}�Wϻ�Ӆ��V]ǻN�����'�6�&�n�w�}�%���¹��_9��R�� ���m�%�u�h�u�� ���Yۖ��V��C1�����d�
�a�h�6�����&����uO��[��W���_�u�u�4�0�l��������l ��]�����h�w�w�"�2�}����
����9��h[�*��h�4�
�:�$��ہ�PӃ��VF�UךU���4�2�g�4�;�2��������l��S��D���=�;�}�
�2�(��������9��S�����;�!�9�f�`�}����[����9F�C����:�0�4�&�0�}����
���l�N��*���0�4�&�2��/���	����@��G1�����u�%�&�2�4�8�(���
�ד�@��N��*���u�%�&�2�4�8�(���
�ӓ�@��d��Uʷ�2�;�u�u�w�}����Qۈ��N��h�����:�<�
�u�w�-��������]�V�����
�:�<�
�w�}��������B9��h��*���
�|�u�'��<�(���
����T��N�����0�u�;�u�6�����&����P9��
N��*���
�&�$���)�(���&���F��R ��U���u�u�u�u�6�����E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���1�;�u�h�6�����&����P9��=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�%�<�;�}����Ӗ��P��N����u�%�<�9��.����	����	F��X��´�
�!�'�y�6�����
����g9��1����_�u�u�0�>�W�W���Y�ƥ�N��X�����:�&�
�:�>��W���	����A���U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�t����Y���F�N��U���<�9�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��RN�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�V�����u�&�<�;�'�2����Y��ƹF��G1�����4�&�2�
�%�>�MϮ�������T����<�
�&�$���ځ�
����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������O�C��U���u�u�u�u�w�<�(��������T�����2�6�d�_�w�}�W������F�N��U���4�
�0�1�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߊu�u�%�'�#�/�(���Dӕ��^9��C1�����0�4�&�2��<����&����l��=N��U���'�!�'�
�w�`����&����e9��^�����2�
�
�4�#�;�(��J����9F������'�
�u�h�$�9�(���&����Z��V�����
�4�!�3��k�N���B�����E�����u�h�;�"�2�o�N���
����lW��1��N�ߊu�u�x�4��4�(���&����R��P �����&�{�x�_�w�}��������lW��h�����%�:�u�u�%�>����	����U��=N��U���<�_�u�u�w�}�W���Y�ƭ�l��h��*��u�h�}�%�4�3����H�����t=�����u�:�;�:�d�t�}���Y����C��R���ߊu�u�x�4��4�(���&����@��YN�����&�u�x�u�w�<�(���&����U��D�����:�u�u�'�4�.�_���:����^OǻN�����_�u�u�u�w�}�W���Y����Z��S
��F��u�4�
��1�0�GϺ�����O������!�9�d�d�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���Y����T��E�����x�_�u�u�'�.��������R��P �����o�%�:�0�$�<�(������F�U�����u�u�u�u�w�}�WϿ�&����Q��V��H���%�6�;�!�;�l�F������l ��_�����:�d�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��A���
������T��[���_�u�u�%�$�:����N�ד�@��Y1�����u�'�6�&��-�4���
��ƹF��R	�����u�u�u�u�w�}�W���
����W��_��H���%�6�;�!�;�l�F������l ��Z�����:�a�|�_�w�}��������@]Ǒ=N��U���4�
�<�
�3��AϿ�
����C��R��U���u�u�4�
�>�����O����Z��G��U���'�6�&�}�'��(���P�����^ ךU���u�u�u�u�w�}��������l_��S�����:�&�
�#��}�W���:����^N��S�����|�n�u�u�2�9��������9l�N�U���&�2�6�0��	����������^	�����0�&�u�x�w�}��������V��c1��D���8�e�4�&�0�����CӖ��P�������7�1�g�|�w�}�������F���]���&�2�7�1�e�t����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����l ��h^��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�o����HӇ��Z��G�����u�x�u�u�6�����
����g9��1�����4�&�2�
�%�>�MϮ�������D�����`�|�u�u�5�:����Y����������7�1�`�|�#�8�W���Y���F������6�0�
��$�o����H���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�&�2�6�2��#���K����lW�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����D�����
��&�f�1�0�EϿ�
����C��R��U���u�u�4�
�>�����*���� 9��Z1�����2�
�'�6�m�-����
ۇ��@��U
��L���u�u�7�2�9�}�W���Yӏ����D�����l�|�!�0�w�}�W���Y�����D�����
��&�f�1�0�E��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�D������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�a�3�8�d�<����Y����V��C�U���4�
�<�
�$�,�$���ǹ��^9��V�����'�6�o�%�8�8�ǿ�&����Q��\����u�0�<�_�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y����C9��P1������&�a�3�:�n�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�i����J���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���`�3�8�a�6�.��������@H�d��Uʴ�
�<�
�&�&��(���&����9��D��*���6�o�%�:�2�.��������W9��GךU���0�<�_�u�w�}�W���Q����Z��S
��C���!�0�u�u�w�}�W���YӇ��@��T��*���&�`�3�8�c�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����0�
��&�b�;���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�u�w�?����>�փ�G9��1��*���
�g�i�u�#�-�N�������F��EN��*���&�
�#�
�~�W�W�������t#��B��Cڊ� �`�b�%�w�`�_���&�ғ�V��Z����4�
�:�&��+�(���s���Q	��h�����
�c�
� �b�o����D�ι�G9��P1�A���:�u�%�6�9�)����H��ƹF��E����
�d�3�
�d�m����D�μ�]	��1��*���d�f�
�g�8�}��������lV��X��D���
�f�m�%�~�W�W�������VU��^\�� ��b�
�g�i�w�-����A����U��X�����'�;�"�<�9�4�(߁�����l ��Z�*��n�u�u�7�:�/��������T��h�I���%�;�!�m�>�;�(��L����\��R�����!�e�;�!�>�;�(��@����l�N�����0�e�1�8�%�<�(�������9��R��]���&�2�7�!�f�/���A�ƭ�WF��[�����0�
�
� �a�i����s���Q��E	��E���8�'�4�
��(�E���	���N��@�����
�0�
�m�g�<�Ϻ�����l	��D1��*��
�f�n�u�w�?�����֓�l ��^�����h�}�'�0�0�i�(�������l��B1�L���u�:�u�%�4�3����H���9F������a�3�
�g�b�-�W��Q����U
��h\�� ��m�
�g�:�w�3��������]	��Q��G���%�|�_�u�w�/����L����U��h�I���:�0�3�:�����K����	��B �����"�f�;�!�1��D���	����F�U�����
� �d�l��o�K�������_	��1��*��c�%�u�'�"�9�����ғ�\��B1�L؊�g�n�u�u�5�0��������9��R��]���d�3�
�g��o��������VR��S�����
�
� �g�n�-�^�ԜY�Ʈ�^��R1��*���c�d�%�u�j�u��������lW��R	��M���:�u�
�:��l����Mƹ��]ǻN�����2�
�g�3��l�F���Y���]��^	�����
� �d�a��n����&����ZT��B1�Cߊ�g�n�u�u�5�0��������lW��1��U��}�0�&�2�5�)�D���&����l��X��*���
�f�3�
�d�i����s���Q��E	��ފ� �d�a�
�e�a�Wǰ�����Q��1��*��e�%�u�'�'�3����&����U��G\����u�'�0�2�����A����[�Y�����<�
�0�
�o�m����&����Z9��h\�*��n�u�u�7�:�/����¹��lP��h�I��� �1�'�9� �l����Aǹ��	��X�����
�
� �c�f�-�^�ԜY�Ʈ�^��R1��؊� �d�d�
�e�a�Wǫ�����\��h��D��
�g�:�u�!�/����K����W��h�N���u�7�8�'�2�4�܁�����9��R��]���0�3�:�
��(�F��&����AF��R�����
� �d�g��o�L���Yӄ��V��h��A���
�a�c�%�w�`�_�������D9��Q��A���%�u�'�:�2�;����&����S��G\����u�'�0�2���(���J�Г�F�F�����9�"�3�
�f��Eϱ�Y����U
��h��G���%�|�_�u�w�<����&����R��N�U¡�%�f�
�0��e�CϿ�Ӓ��lW��E��D��|�_�u�u�6�/�(���K�Փ�F�F�����!�'�2�d�n�}��������A��V�\�ߊu�u�0�0�2�����H����U��G]��H�ߊu�u�u�u��l��������F��R �����,�d�3�
�e��E��Y���O��[�����u�u�u�4�0�l��������A��V�N���u�1�9�!�3�2��������l��S��U���u�u�!�%�d�;�(��&����[������� �g�f�%��t�J���^�Ʃ�@�N��U���&�2�7�!�%�:�F��B�����R��*���:�
� �c�o�-�W��s���F�e��ۊ�9�
�;�&�%�:�F��Y����N��E��D���
�g�
�g�g�}�W��PӃ��VFǻN��U���4�2�d�4�;�'��������
V��=N��U���
��-� ��k�(�������l��S�����:�<�
�0�#�/��������R��X ��*���g�e�u�u�9�4��������C��1��\�ߊu�u�-�
��%����Oʹ��9��h]�*��i�u�u�u�w�}����8����F��W��*ي� �f�a�%�w�5��������U�� ^��G��u�u�d�|�2�.�W���Y��� ��h/�����
�c�
�
�"�n�A���B��� ��h/�����
�c�
�
��(�D���	���l�N��Uʥ��9�
�l�:�%����Mù����YN�����2�
� �f�c�-�_���D����F��D��U���u�u�%��;��(�������9��d��Uʳ�%����#�l�N�������9��R�����9�2�6�#�4�2�_���������T�����f�
�|�x�"�.����Q����r$��x��D����f�3�
�b��D���s���U��y+��:���d�`��3��m�(��E�ƿ�W9��P�����:�}�;�<�9�9��������_��h^��Xʠ�&�2�0�}�/���������V��a1��*��
�d�|�_�w�}����<����G9�� 1�����l�
�g�i�w�)�(�������P�������1�4�
�:�$�����I���F��P ��]���
�:�0�!�%��Oہ�&����
W��G����u�-�
�!��.�(�������V9��h8��*���d�m�
�f�k�}�W���Y����K��C1�����!� �!�'��k�!�������
Q��@��U¦�9�!�%�
�2��N��I���W����ߊu�u�u�u�/�����
����A��B��A؊�
� �d�b��n�}���Y����P��V��&���6� �0�a���(���H����CU�
NךU���u�u�-�
�#���������F��W��*݊� �d�g�
�d�*����
����^��h��*��`�e�u�u�f�t����Y���F���*����&�
�!�"�)����K����l ��[�*��_�u�u�u�w�%�(���:����`��T����
�
�
� �f�d�(��E�ƿ�W9��P�����:�}�0�<�2�.����Q����U��R	��L��y�g�|�_�w�}��������@��C�����
�g��m�1��B���	���l�N��Uʳ�%�6�
�4�2���������9�� 1��*��b�%�u�=�9�u��������A��W�]���h�r�r�u�;�8�}���Y���U��T������'�6� �2�i�(���&����_��G]�U���3�%�6�
�6�8�$�������lR��a1��*���b�%�u�h�]�}�W���Y����P��V��&���6� �0�a���(���H����CW��_��]���6�;�d�g��8�(��H���F�G�����_�u�u�u�w�����K�֓�K��d;��:����7�
� �f�n�(��s���U��T������'�6� �2�i�(���&����S��G]��H�ߊu�u�u�u�/�����
����A��B��A؊�
�
� �d�n��Fϩ�����V
��Z�����d�a�}�|�j�z�P������F�N�����6�
�4�0��/��������e9��h_�B���n�u�u�3�'�>�(�������F��E��L���a�3�
�`�f�-�W��s���F�Q�����4�0��'�4�(���&����A��W�U���;�}�0�
�:�l�(���&����V�
N��R���9�0�_�u�w�}�W���&����R��d�����0�a�
�
��(�F��&����F�Q�����4�0��'�4�(���&����U��\�����h�_�u�u�w�}�(���K����l��h��D��
�f�"�0�w�?����Ź��lW��1��]���h�r�r�u�;�8�}���Y���C9��[\��*���3�
�`�g�'�f�W�������G9��D�����!�'�
�l��e����L�ѓ� F�d��U���u�3�%�6��<��������A��1��B���2�d�b�u�?�3�_���&���� 9��P1�C���|�h�r�r�w�1��ԜY���F��G1��*���0��'�6�"�8�Cց�&ǹ��lW��1��N���u�3�%�6��<��������A��1�����`�b�%�u�j�W�W���Y�ƪ�C9��h-�����'�6� �0�c��(؁�����9�������'�6�;�d�e�����@���F�_��U���0�_�u�u�w�}����*����F��B�����d�c��&�1��B���	��ƹF��O�����&�
�!� �#�/�(���/�ԓ�F9��Z��F��u�u�u�u�w�;����&����l5��B�����l��b�3��h�G���Y����N��[1��Ҋ�0�
�l�m�g�}�W��PӃ��VFǻN��U���-�
�!��$���������P��h��D��
�f�_�u�w�%�(���:����`��T�����
�
�
� �f�o�(��E��ƹF�N�����!��&�
�#�(����&�ԓ�lQ��B1�L݊�d�"�0�u�$�1����H����lW��F�U���d�|�0�&�w�}�W���YӀ��l��t��*��� �!�'�
�a��E���&����l��=N��U���
�!��&��)��������l0��h��D��
�f�i�u�w�}�W���	����9��1�����
�f�e�%�w�5��������VS��B1�Cފ�g�e�u�u�f�t����Y���F������f�g�
� �f�j�(��s���U��T������'�6� �2�h�(���&����T��G]��H�ߊu�u�u�u�/�����
����A��B��Aӊ�
�
� �d�e��Dϩ�����V
��Z�*���
�l�g�e�w�}�F�������9F�N��U���
�!��&��)��������l0��h��D��
�f�_�u�w�%�(���:����`��T�����
�
� �d�g��D��Y���F���*����&�
�!�"�)����O����l��h_�Aʢ�0�u�:�
�8�9�(�������
R��G��U��|�0�&�u�w�}�W���	����9��1��؊�
� �d�a��n�}���Y���U��Y��*���8�f�a��1��Nށ�H���@��[�����6�:�}�0�>�8�����Υ�l��_��*���f�|�n�_�w�}�W�������W��R��A����3�
�l��l�K�������T��A�����0�<�0�&�0�8�_���&����|��X��#���3�
�`�
�d�q�D���s���F���*���0�!�'�
�b��(�������U��G_��Hʦ�1�9�2�6�!�>����������Y�����;�1�
�0�:�i�O�������
9��B�\��_�u�u�-��2��������9��Q��Gӊ�f�i�u�!�'�l�(���N�ד� F�V�����
�#�f�e�l�}�Wϸ�	����q��C1�����6�
�l�
�����K˹��Z�=N��U���u�-�
�!��.�(�������V9��h8��*���d�g�
�f� �8�WǪ�	�ѓ�V��_�E���u�d�|�0�$�}�W���Y����K��C1�����!� �!�'��o�!�������
Q��UךU���6�%�`�;�#�;�(��J����[�^��D���
�e�`�%�w�2�W�������l
��h_����u�6�%�
�"�l�Bځ�K���V�@��U¡�%�`�
� �f�i�(��DӇ��P	��C1��G��u�9�0�w�u�W�W�������U��Z�����h�w�w�"�2�}�����θ�C9��h��D��
�a�u�u�>�3�ǿ�&����G9��1�\ʰ�&�u�e�n�w�}����J����P��h�I���d�u�=�;��4��������9��h_�F���|�i�&�2�2�u��������ER��G�����w�w�_�u�w�>�ہ�����9��R��W���"�0�u�&�0�8�_���&�ԓ�F9��Y��A���u�<�;�1�6�����&����O�R��U��n�u�u�<�:����L����[�L�����}�8�
�`�1��@؁�J����C9��Y�����e�u�9�0�u��}���Y����l��h��B���%�u�h�}�4�-����Aƹ���������!�9�d�d�l�}�WϷ�����l ��\�*��i�u�
�4�e�n�(���H����CT�N�����u�f�n�u�w�4����K����R��h�I���
�4�g�a��(�F��&��� F��@ ��U��n�u�u�<�9�:����H�ߓ� F������f�
� �d�d��E��Y����G	�G�U���;�2�&�6�1��@ց�K�����Y��*���
�b�`�4�3�3� �������A��V�\�ߊu�u�0�
�%���������l��S�����&�6�3�
�`��EϦ�Ӈ��P	��C1��D��n�u�u�;� �8�F߁�����l��S��U���u�u�<�
�;�5�(ށ�Y����N��[1��ߊ� �m�b�%��t�J���^�Ʃ�@�N��U���3�%����)�F���/�Փ�V��]����u�0��9�f�;�(��&���FǻN��U���-�
�:�0�#�/�(��&����lS��h����u�&�9�!�'����H����O�I�\ʰ�&�u�u�u�w�}����7����F��Y��*���`�a�%�n�w�}��������U��X��F��u�u�u�u�w�;����>����lW��h8�� ���a�%�u�=�9�u��������9��^��H��r�u�9�0�]�}�W���Y����}#��x��D����'�2�d�b�f�W�������_W��Q��@ي�f�i�u�u�w�}�Wϰ�����W��V�����f�
�d�"�2�}��������F9��1��]���h�r�r�u�;�8�}���Y���]��R�*���l�m�%�n�w�}��������U�� Y��F��u�u�u�u�w�<�(���
���� 9��@��U¦�9�!�%�
�"�j�F���Q���A��N�����u�u�u�u�6�����&����]ǻN�����9�`�3�
�o��D��Y���F������!�9�f�`� �8�WǷ�����lS��h�E���u�d�|�0�$�}�W���Y����C9��Y�����a�_�u�u�2��������� 9��R�����u�u�u�0��1�Eށ�����R��Q��Cӊ�f�"�0�u�8���������
9��^��H��r�u�9�0�]�}�W���Y����V
��h��L���%�n�u�u�9�*��������9��R�����u�u�u�-������&����e9��P1�@���=�;�}�0��0�@���&����CT�N��R��u�9�0�_�w�}�W�������W��R��A����'�2�d�b�f�W���Y����V��[\�*���!�3�
�d��l�K�������T��A�����0�<�0�&�0�8�_���*����U��^��F���f�|�_�u�w�}�Wϰ�����W��V�����f�
�d�i�w�)�(�������P�������&�2�0�}�2���������9��B�\��_�u�u�0��1�Eށ�����R��Q��Cӊ�f�i�u�u�w�}�WϿ�&����G9��1����u�&�9�!�'����N����O�I�\ʰ�&�u�u�u�w�}��������_��UךU���0��9�g��<����&����l��S�����:�<�
�0�#�/�����ι�@��R
�� ���0�!�'�d��/����
����l��h_�E���|�n�u�u�9�*��������9��R�����u�u�u�-������&����e9��P1�@���=�;�}�6�'�;�(��&���F�_��U���0�_�u�u�w�}��������V��^��#���2�d�`�n�w�}�����Փ�F9��1��U��_�u�u�u�w�8�$������� 9�������'�6�;�
�"�e�N���Q���A��N�����u�u�u�u�9�*��������9��d��Uʻ�"�0�a�3��m�(��E��ƹF�N�����:�0�!�'��h�(�������F9�� 1��U���;�}�0�
�:�h����IĹ��V�
N��R���9�0�_�u�w�}�W���&����|��X��#���'�2�d�f�l�}�Wϰ�����l ��X�����h�_�u�u�w�}��������V��^��#���2�d�`�u�?�3�_���&����l ��^�����|�h�r�r�w�1��ԜY���F��G1��2���!�d�b��1��Nہ�K���F��@=��C���
�b�
�f�k�}�W���Y����K��r)�� ���f�
�
�0��e�Oϩ�����V
��Z�����b�
�g�e�w�}�F�������9F�N��U���
�:�0�!�%��Oہ�&����
W��UךU���0��9�
�"�e�N���Y���F�N�����;�1�
�0�:�n�C�������9�������6�%�3�
�o��E��Y���O��[�����u�u�u�-������&����e9��h[�*��_�u�u�0��1�(���A�ѓ� F�d��U���u�;�"�0�b�;�(��&����[�������
� �m�l�'�u�^��^���V
��d��U���u�;�"�0�a�;�(��&����F�Y�����3�
�d�
�d�a�W���Y�����d��*���l�f�%�u�?�3�_�������U��W��G��u�u�d�|�2�.�W���Y��� ��h/�����
�c�
�
��8�(��J���F��@=��*���m�f�%�u�j�W�W���Y�ƪ�C9��S�����a�`��'�0�l�B������@��C��*���m�b�%�}�~�`�P���Y����l�N��Uʳ�%����#�l�B�������S��=N��U���&�2�7�!�g�3����&���� T��G\��H���0�&�2�7�#�n����K�Г� F��EN��*���&�
�#�
�~�W�W�������]��h^�����g�3�
�a�e�-�W��Q����Z��^��*���d�g�
�f�/�/��������_��G�U���;�"�<�;�>��(���&����lW��1��U��}�0�&�2�5�)�E���&����l��O�����:�&�
�#��t�}���Y����Z��^��*���a�e�%�u�j�-�!���&�Փ�F9��1��]���1�"�!�u�b�f�W�������T��C1�����d�b�%�u�j�-�!���&�֓�F9��]��G��u�:�;�:�d�t�}���Y����Z��^��*���d�m�
�f�k�}�(���K����U��X�����d�1�"�!�w�l�L���Yӈ��@��U��A���
�a�e�%�w�`��������l ��Z�*��f�u�:�;�8�n�^�ԜY�Ƣ�D��Y��*���g�d�%�u�j�-�!���&����lT��h�F���:�;�:�f�~�W�W���	����V��V����� �g�`�%�w�`�}���Y���Z��[��*ۊ�u�=�;�}�:����J����O�I�\ʰ�&�u�u�u�w�}����8����F��Y��*���g�l�%�n�w�}��������T��B1�Cۊ�g�i�u�<�:�l����I�ӓ�F��SN�����
�e�
�g�l�}�Wϱ�&����9��hV�*��i�u�&�9�#�-�(���N�ד�F����*���g�3�
�a��o�L���YӉ��P	��1��*���
�g�i�u�8���������
9�������:�1�
� �o�l����s���\��X �����d�
�g�i�w�.����	ƹ��l^��h����0�
�8�f�1��Oց�K��ƹF��B�����'�d�
�'�#���������V��h�I���u�u�u�u�9�*���&����
U��N�����:�
�:�1��(�O���	����[�I�����u�u�u�u�w�3� ���Hƹ��l_��h����u�#�'�9� �l����O¹��Z������
�d�3�
�b��EϿ�Ӓ��lW��Q��@܊�g�n�u�u�8�8����&����lW��1��U��}�'�0�2��o����H�ד�F��SN����
� �d�b��o�L���YӉ��A ��@1�����f�g�%�u�j�u��������l ��]�*��4�1�!�%�e����HŹ��]ǻN�����9�"�a�3��i�A���Y���Q��E	��ފ� �d�a�
�e�<�Ϫ�	����U��[�����_�u�u�#�%�1� ���&����CT�
N�����2�
�
� �e�e�����Ƹ�C9��Q��C݊�g�n�u�u�'�m�@܁�&����lR��B1�Cي�f�i�u�u�w�}�WϿ�&����G9��_��U���;�}�8�
�n�;�(��L����O�I�\ʰ�&�u�u�u�w�}����Lƹ��lW��1��N���u�%�e�b���O���M����Q��h�I���u�u�u�u�6�����&����lV��_��]���
�d�3�
�a�d����P���A�R��U���u�u�u�!�'�h�(���H����CW��N����b�
�
�m�a�i����N�ד� F�d��U���u�4�
�:�$�����Iӑ��]F��Z��F���
�b�f�%��t�J���^�Ʃ�@�N��U���!�%�`�
�"�l�Dځ�H���F��V��*���c�e�%�u�j�u����&¹��lP��h�����;�0�
�;���������_��d��Uʥ�a�
�
� �b�k����D�Ξ�]��h��*���&�3�
�d��o��������9��h[�*��n�u�u�%��.����&����^��N�U���
��-� ��n�(�������l��\�����:�g�|�_�w�}�(�������l ��_�*��i�u�
�4�e�n�(���H����CT�N�����u�g�n�u�w�-�%�������U��\��A��u�-�
��/�(�(��&����lR��h�F���:�;�:�f�~�W�W���&����lW��Q��Dފ�a�i�u�-������&����e9��hZ�*��g�u�:�;�8�l�^�ԜY�Ƽ�e��h_�*���
� �b�b�'�}�J�ԜY���F��h�����#�c�b��w�5��������V9��^_�� ��l�%�}�|�j�z�P������F�N�����9�
�f�'�0�l�@��Y����l0��1��Dӊ� �b�a�%�w�`�}���Y���R��X ��*���c�m�e�u�?�3�_�������D9��Q��Mފ�g�e�u�u�f�t����Y���F������g�
�0�
�o�d�}���Y����_T��h��D���%�u�h�%��1�(�������l��X�����:�d�|�_�w�}�(���K����l��h��D��
�f�i�u�w�}�W�������]��[�*ݓ����"�2�}��������l��Q��F���%�}�|�h�p�z�W������F�N��#���
�a�3�
�e�o���Y����l0��1�C���-�3�
�`�c�-�W��s���F�V�����
�#�g�b���1������Q��E	�����
� �d�m��o�G���Y�����RNךU���u�u�
�4�e�i�(���H����CW��N�����9�
�g�
�6�o����&����l��S��U���u�u�3�%�4�����*����G��hZ��#���3�
�f�b�'�}����Q����9��P1�D���|�h�r�r�w�1��ԜY���F��G1��*���0��'�6�"�8�Bف�&Ĺ��T9�� Z�U���%��9�
�d�����*����F��B�����`�`�%�u�j�W�W���Y�ƪ�C9��h-�����'�6� �0�b��(؁�����R��_��]���
�
�0�
�n�n�G���Y�����RNךU���u�u�-�
�#���������F��W��*݊� �d�g�
�d�W�W���&����lT��Q��Bފ�g�i�u�!��2����������^	��¥��9�
�m�1��Fہ�M���F��P ��]���
�
� �a�g�-�^��Y����l0��1�*���m�b�%�u�j�W�W���Y�Ƣ�D5��1��*��
�f�"�0�w�2�(�������l^��h�E���u�d�|�0�$�}�W���Y����V��[\�� ��b�%�n�u�w�-�!���&�ޓ�F9��_��G��u�!�
�:�>�����ە��]��E1�����e�b�%�|�|�.����Q����_��B1�F݊�d�|�_�u�w�����K����W��G\��Hʦ�1�9�2�6�!�>��������V��h8��G���3�
�c�
�c�}�W���������h_�� ��d�%�|�n�w�}��������l ��_�*��i�u�!�
�8�4�(�������Z��SF����
� �d�g��l�W���������h\�����d�e�%�|�l�}�WϮ�/���� U��B1�Cӊ�g�i�u�!��2����������Y�����a�
�4�!�1��E���	�����Y�����'�2�d�g�~�f�W���	����9��h��D��
�d�i�u��<�E��&����P��G\��G���d�1�"�!�w�t�}���Y����_T��1�����
�a�
�f�k�}�W���Y����C9��Y����
�����*��������T��h�� ��c�%�}�|�j�z�P������F�N�����9�
�
�0��e�C�ԜY�Ƽ�e��h]��E���
�f�m�%�w�`�}���Y���R��X ��*���g�m�e�e�g�}����Q����A ��@1�����f�c�%�}�~�`�P���Y����l�N��Uʥ��9�
�a�1��E���	��ƹF��h8��G���3�
�l�
�d�a�W���Y�����d��*���m�b�%�u�?�3�_�������l ��[�����|�h�r�r�w�1��ԜY���F��@=��B���
�b�
�f�]�}�W����ԓ�9��h_�F���u�h�&�1�;�:��������@��R
�����`�6�&�
�"�l�G߁�H���@��R
��*���
�0�
�l�g�t�}���Y����_T��1��*��c�%�u�h�'��݁�H����R��h�F���u�u�:�;�8�m�L���YӖ��R
��1�*���d�d�
�f�k�}�W���Y����C9��Y����
�e�e�e�g�*��������U
��hZ�� ��m�
�g�e�w�}�F�������9F�N��U���4�g�a�
�"�l�Fف�H���F��a��*ފ� �l�d�%�w�`�}���Y���]��R�B���&�
� �l�`�-�W����Σ�l��S\�� ��d�%�}�|�j�z�P������F�N��������!�f�h�!�������]ǻN��*���g�`�3�
�a��D��Y���F� ��&���f�3�
�`��n� ���Yۉ��P	��1��*���
�g�e�u�w�l�^ϻ�
��ƹF�N�����9�g�3�
�c��D�ԜY�Ƽ�e��h��M���
�a�
�f�k�}�W���Y����C9��Y����
�e�e�e�g�*��������U
��h��F���%�}�|�h�p�z�W������F�N��#���
�
�0�
�o�i�}���Y����_T��h��D���%�u�h�<��8����/���F��a��*��� �d�`�%�w�`��������l��C�����/�}�;�<�9�9��������l��C�����0�}�
�4�e�.����Mƹ��F�D�����e�u�4�
�8�.�(���N����O�N�\��u�u�%�;�#�e�ށ�����9��R��W���"�0�u�!�'�l�(���H����CR������!�9�g�f�w�1����[���F��Y��M���
� �d�c��o�K���I�ƻ�V�C��Gߊ� �d�g�
�c�`��������_��G�����w�w�_�u�w����&����lW��1��U��w�w�"�0�w�-�%�������U��[�����u�%�6�;�#�1�D��Y����D��d��Uʥ�;�!�<�
�"�k�B���Y���W��C�����&�3�
�g��n��������]��[��D��u�u�%�;�#�4�(���H����CT�
N��Wʢ�0�u�%��$�1�(܁�����9��S�����;�!�9�f�g�}����[����F�G1�����
� �d�e��o�K���I�ƻ�V�C��Dڊ� �d�l�
�c�`��������_��G�����w�w�_�u�w�����M����R��h�I���e�u�=�;��0�(�������^��N�����:�&�
�#��t����Y���9F������
� �g�f�'�}�J�������G9��P1�L���:�u�4�'��(�E���	����F�F�����;�d�3�
�g��E��Y۔��l��B1�L���u�;�u�7�#�;�(��&���9F������2�
�
� �c�i����D�ξ�Z9��h��A���%�u�;�u�5�)�F���&����CU�=N��U���!�d�3�
�e��D��Y����}#��x��D����3�
�e��o�F�������W��d��Uʤ�<�
� �d�d�-�W��	����9��Q��Aߊ�g�d�u�:�9�2�F���s���A9��Q��F܊�g�i�u�e�w�5��������l ��]�����u�%�6�;�#�1�F݁�PӃ��VF�UךU���
�
�
� �f�n�(��E�ƿ�W9��P�����:�}�<�;�3�)���&����T��G_��^ʦ�2�0�}�8��e����I�ѓ�O�=N��U���
� �d�d��o�K�������T��A�����<�;�1�!�'�l�(���H����CW�N�����}�8�
�c�1��G���	���9F��� ��`�%�u�h�u�� ���Yے��lU��Q��Mۊ�d�h�4�
�8�.�(���M���V
��L�N���u�'�<�<��(�C���	���N��G1�*���a�e�%�u�%�/�F���&����CT�=N��U���
�
� �d�n�-�W��Q���� T��B1�D���u�'�'�3��e�(��B�����h��C���%�u�h�}�8�1����6����R��B1�G���u�:�u�%�4�3����H���9F���*���d�
� �d�n��E��Yە��l��]�����'�4�
� �f�d�(������C9��Y�����d�n�u�u�$�1����H����W��h�I���!�%�`�3��m�(������V
��Z�*���d�l�
�g�l�}�Wϭ�����T��B1�Dߊ�g�i�u�&�;�)���&����A��h��D��
�g�-�'�6�����&����O��N�����!�%�f�
�2�2��������
W��N�Uº�
�:�1�
�e�;�(��H����\��Z��B���
�e�b�%�~�W�W�������CW��S�����
� �b�b�'�}�J�������CP��R�����3�
�`�
�e�2�W���&ƹ��lP��h�N���u�&�9�!�'�n����H�ד�F�F�����3�
�d�
�e�<�ϭ�����T��B1�Dߊ�g�n�u�u�$�1����Mǹ��^	��V �� ��e�
�g�i�w�.����	����W��E	��*���d�l�
�g�8�}����&����P��G�U���&�9�!�%��(�@���	���N��Z�� ���`�%�u�:�w�-��������lW�=N��U���
�8�g�
�2�2��������9��R��]���
�8�d�
�2�2��������9�������c�3�
�d��o�L���Yӕ��l��1��*��
�g�i�u�%�+����Iù������*���d�3�
�a��o�L���Yӕ��l��1��*��
�g�i�u�#�-�A���&����CT��Y
�����8�
� �b�d�-�^�ԜY�ƿ�_9��GZ�� ��d�%�u�h��8�(���K����^	��V �� ��`�%�u�:�w�-��������lW�=N��U���
�8�`�3��m�(��E����^��h��C���%�u�;�u�2���������9��UךU���0�
�8�c�3�0����&����U��N�U¼�8�
� �`�b�-�W�������F9��1��\�ߊu�u�0�
�:�k����Oƹ��Z��������!�d�c�;�(��&����]��T�����3�
�`�
�e�f�W���
����^��Q��Bۊ�g�i�u�!�'�h����IŹ������*���c�3�
�c��o�L���Yӕ��l��1��*��`�%�u�h��0�(�������Q��N��ʦ�9�!�%�
�"�l�@ց�K��ƹF��R�����3�
�e�l�'�}�J�������t#��B��Cފ� �`�g�%�w�/����Hƹ��G9��h_�F���|�_�u�u�2���������l��S�����!�%�f�1�:�/��������l��O�����:�&�
�#��t�}���Y����l��h8�����
�&�<�;�f�;�(��L����[�N��U���%�e�b�
��e�O�������Q��N�����<�8�f�3��k�D���Q���A��N�����u�u�u�u�6�����&����lW��^�E�ߊu�u�&�8�>�)�!�������@��Y1�����
� �d�g��l�K�������T��A�����0�<�0� �$�:����
����]��h�����&�<�;�d�1��@���	���O�=N��U���8�<�!�� �4����
����9��h_�L���u�h�_�u�w�}�W���K�Փ�lV��1�����b�d�%�u�?�3�_���	ǹ��lW�� 1��]���h�r�r�u�;�8�}���Y���R��X ��*���d�d�e�e�g�f�W���
����Z��a1�����4�&�2�
��<����&����l��S�����:�<�
�0�#�/�����ι�@��R
�����<�!��"�>�8��������lW��1��\��|�n�u�u�$�9�(���&����Z��V�����4�!�3�
�`�j����Dӕ��l
��^�����'�'�&�/��3����ە��^9��C1�����0�4�&�2�����Lʹ��J��G�U���&�1�
�;������&����T��B1�Bۊ�f�i�u�u�w�}�WϮ�I����9��V��*���d�c�
�f� �8�WǷ��ԓ�F9��W��G��u�u�d�|�2�.�W���Y�����T�����f�
�e�e�g�m�}���Y����U��R�����3�
�b�
�e�a�WǮ�J˹��U��^��Gʺ�u�'�0�2�c���������9��hX�*��n�u�u�!�'����A����[�X�����
� �g�f�'�}�ϰ�����l��h��F���%�|�_�u�w�0�E���&����CT�
N����f�1�8�'�6����K����K	��V�����
�#�
�|�]�}�W���J����_��G\��H���'�0�2�a��8��������U��Y��Gʺ�u�8�
�f�1��Bف�K��ƹF��Z��E���
�g�a�%�w�`��������l ��\�*��f�u�:�;�8�n�^�ԜY�Ƹ�C9��h��A���%�u�h�}�2�.�����ד�F9��1��U���u�%�6�;�#�1�F��B�����h_�����a�
�g�i�w�)���&����
R��N��ʴ�
�:�&�
�!��^�ԜY�Ƹ�C9��h��C���%�u�h�}�>�3����&����^����U���6�;�!�9�f�l�L���YӒ��lW��Q��Gۊ�f�i�u�u�w�}�WϮ�/����_��Z�����e�
�f�"�2�}��������lW��X�� ��d�%�}�|�j�z�P������F�N�����9�
�
�l�1��Fہ�J���F�N����
� �d�e��l�K�������T��A�����0�<�0�&�0�8�_����ԓ�l ��X�����f�|�n�_�w�}�W�������l ��^�*��i�u�!�
�8�4�(�������V��RF�����}�
�4�g�c�;�(��&��� R�dךU���u�u�8�
�`�;�(��J����[��C
�����
�0�!�'�%�.����������V��F���
�l�
�f�{�i�^�ԶY���F��Z��M���
�e�b�%�w�`��������l��C�����/�}�<�;�3�-�!���&�Г�F9�� 1��\��|�n�_�u�w�}�W���&�ߓ�F9��Y��D��u�!�
�:�>�����۔��Z��D�����;�8�-�g��q�C���s�����h_�� ��d�%�u�h�$�9��������G	��E�����;�<�;�1�&������ד�F9��1��\��|�n�u�u�w�}����Kù��lW�� 1��U��&�1�9�2�4�+����Q����I��^	��¥��9�
�m�%�:�F��P����]ǑN��U���!�%�g�
�"�l�D߁�H���@��[�����6�:�}�0�>�8�����ξ�e9��E��D��|�f�|�n�]�}�W���&�ԓ�F9�� Y��G��u�<�;�2�1��F���	�ƴ�AF��h�����#�
�|�_�w�}����J����T��h�I���u�u�u�u�#�-�Cف�����9�������'�0�2�a�1��E���	����[�I�����u�u�u�u�w�)���&����R��G]�U���!�%�g�
�"�l�Fف�K�����R	��*���d�b�
�f�/�/��������_��G�U���!�%�g�
�"�l�Eׁ�M���C9��[\��D���
�a�f�%��n��������]ǻN�����c�3�
�a�g�-�W��Q����T9��Q��A���%�u�:�u�'�>�����ד�]ǻN�����b�3�
�e�`�-�W��[����[����*ފ� �`�b�%�w�}��������EU��N�����e�n�u�u�#�-�E���&����CT�
N�����2�7�!�3��o�(������C9��Y�����d�n�u�u�#�-�D߁�����l��S��*���g�&�3�
�c��E��Y����W	��C��\�ߊu�u�8�
�e�;�(��&���F��a��*��� �d�`�%��h��������]ǻN�����`�3�
�b��n�K�������K!��x��D���3�
�c�
�e�{����&����|��X�����`�
�g�n�w�}����J˹��lR��h�I���-�
��-�"��Dځ�&����V��F�U���u�:�;�:�g�f�W�������l ��X�����h�}�<�;�>�����N����\��G1�����9�d�d�n�w�}����Mù��lR��h�I���-�
��-�"��Dځ�&����V��F�U���;�:�d�|�]�}�W���&�ԓ�F9��1��U��3�%����)�F���/����V��G\��Lʱ�"�!�u�l�l�}�W���YӒ��lR��T��*���d�c�
�d�k�}��������E��X�����0�&�2�0��0�(�������Q��G�A���_�u�u�u�w�)���&����l ��Z�*��i�u�!�
�8�4�(�������V��RF�����}�-�
�!��.�(�������V9��h8��*���
�l�a�y�c�t�}���YӒ��lR��Q��G���%�u�h�%��1�(������� U��F�U���;�:�d�n�w�}����MŹ��lW��1��U��_�u�u�u�w�-��������9��q(��3���=�;�}�'�2�:�(���K����T��h�E���u�d�|�0�$�}�W���Y����^��1��*��d�%�n�u�w�)���&����R��G]��H�ߊu�u�u�u�'�>��������V��^�U���;�}�;�0�1�2�(݁�����9��^��H��r�u�9�0�]�}�W���Y����S��B1�Fۊ�a�_�u�u�:��(���L�ѓ�F�F�����-���!�f�i����O����@��X������!�d�e�1��B؁�K���Q	��h��E���
�`�
� �b�o����s���G��Z�� ��a�
�f�i�w�?����>����G9��1��*��
�g�s�7�8��0�������9��h[�*��n�u�u�!�'�h�(���H����CW�
N�����
�4�0��%�>����Mʹ��9��h_�B���}�d�x�d�3�*����P���F��G1�*���d�e�
�d�k�}��������V9��E�� ���a�
�
�
�"�l�N؁�J����F��S�����|�_�u�u�:��@���&����l��S�����!��&�
�#�(����&�Г�l^��B1�GҊ�f�f�u�u�w�2����I��ƹF��Z��M���
�c�l�%�w�`��������@��C�����
�l��m�1��B���	������Y��G���_�u�u�8��d����O�ӓ� F���*����&�
�!�"�)����@����l ��[�*��f�u�:�;�8�n�^�ԜY�Ƹ�C9��Q��E܊�g�i�u�d�w�5��������U��Y��A��4�
�:�&��+�(�������V�=N��U���
�e�3�
�a�n����DӀ��l��t��*��� �!�'�
�e��O���&����l��_�����:�g�|�_�w�}����H����P��h�I���-�
�!��$���������T��hV�� ��l�
�f�f�w�2����J����F�C��C؊� �d�g�
�c�a�W���&����R��d�����0�`�
�
��(�F��&���F��@ ��U��n�u�u�!�'�k�(���H����CU�
N�����
�4�0��%�>����LŹ��9��h_�M���}�d�1�"�#�}�F��Y����^��h��C���%�u�h�w�u�*��������l ��X�����u�%�6�;�#�1�D��Y����D��d��Uʡ�%�b�3�
�f��E��Y���D��F�����3�
�c�
�c�`��������_�� G�����w�w�_�u�w�0�(ׁ�����l��S��D���=�;�}�<�9�9����8����F��W��*ي� �f�a�%�~�c�����έ�l��D�����e�|�0�&�w�m�L���YӒ��l ��Z�����h�w�w�"�2�}�����Υ�l��_��*���k�&�2�0��-��������9��N�����e�n�u�u�#�-����&����CW�
N�����2�6�#�6�8�u����ۓ��Z��SF��*���<�;�f�3��k�(��U���l�N�����
�l�
�g�k�}�F������F��P ��]����'�4�
�$�4����&����CU�N�����0�}�-�
��%����Oʹ��9��h]�*��|�0�&�u�g�f�W�������U
��h_�� ��a�%�u�h��4����&¹��T9��V�����8�g�3�
�`��E��Y����]��Q��*ۊ�:�
� �b�f�-�W��Q����l ��W�����'�%�f�
��(�A���	����F�B �����"�g�3�
�e�j����D�ή�^��R]�����
�g�d�%�w�3�W�������lW��1��\�ߊu�u�;�0�1�2�(݁�����lW��1��U��}�;�0�3�8��(���H����CT��X�����;�!�9�d�f�f�W�������U
��h]�� ��a�
�g�i�w�?�����ߓ�9��h_�E���u�;�u�&�2��(���H����CU�=N��U���0�3�:�
��2�(���H����CT�
N�����3�:�
�
�"�l�Cف�KӞ����T�����d�d�n�u�w�(��������l ��Z�*��i�u�7�8�%�8�N���&����Q��G\�����&�0�
�
�"�l�Gׁ�J��ƹF��Y
�����
�
�:�
�"�l�N݁�K�����R�����
� �d�m��o��������]��[��D��u�u� �1�%�1� ���&����CT�
N�����'�
� �g�n�-�W���Y����A��1�����e�
�g�n�2�9������