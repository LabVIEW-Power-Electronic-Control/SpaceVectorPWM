-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��[�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�_�&�w�8��������Z��X����_�0�!�!�w�k�2���:����l ��A1����g�&�f�
�w�.�W�������Z�=N��U���u��u�u�w�}�MϷ�����\�UךU���u�u� �
���W������V�
N����u�u�u�<�g�
�3���Cӏ��V��T��F��u�u�u�u�3�3�(���-����Z��P��O���g�_�u�u�w�}����.����\��Y�����h�f�_�u�w�f�W���	����l�N��Uʶ�>�u�o�<�w�.��������F�N�����!�o�<�u�$�9�������F�N��U���o�<�u�&�3�1����s���F�S��U��<�u�&�1�;�:��������W��h9��!���u�:�;�:�g�f�W���Y����Z��T�����!�
�:�<��8��������d/��C����!�u�|�_�w�}�W������	F��CN�����2�6�#�6�8�u����.����W��X����_�u�u�n�2�9������ƓR��^�����u�'�=�:�w�k�2���:����l ��A1����g�&�f�
�w�.�W���T���K�C�X���x�x�u�:�'�3����T���K�C�X���x�x�u�u�4�0����Ӌ��v#��t+��E���
�1�#�`�9�����Kӏ��F�N�����u�_�u�u�w�}�W������F�N��U���u�u�u�;�w�)�(�����ƹF�N��U���6�>�;�u�w�}�W���Y�������*���<�n�u�u�w�}�W���
����@9��C�����u�u�o�<�w�.��������F�N��U���&�4�<�
��9����Y���	F��N�����2�6�#�6�8�u�FϺ�����O��N��U���u�u�&�4�>��(������F�N��Uʦ�1�9�2�6�]�}�W���Y���@9��^��*���!�u�u�u�w�}��������T��A�����d�1�"�!�w�t�}���Y���F�Z1�����0� �!�!�6�4�W����ƿ�W9��P�����u�u�u�u�w���������G9��V��U��� �u�!�
�8�4�(������F��@ ��U���u�u�u�u�~�W�W����Ư�^��R �����u�x�x�x�z�p�Z��T���F��T�����4�u�x�x�z�p�Z��T���9F������4�9�u�u�w�g��������l�N�����u�6�>�;�w�}�W���&����P]ǻN�����9�4�!�4�>�}�Mϭ�����Z��N�����4�u�
�1�#�}�W�������T��A�����d�1�"�!�w�t�}���Y����R
��h�����u�u�!�
�8�4�L���Yӕ��]��U1�����u�o�&�1�;�:�������� W��X����n�u�u�&�0�<�W�������F��D�����6�_�u�u�>�3�Ϭ�����F���*���<�
�0�!�%�n�W������]ǻN�����9�1�;�
�"�l�Mϭ�����Z��R��±�;�
���z�}�������9F������1�;�
� �f�g��������l��C�����
���x�w�2����I����V��=N��U���x�x�x�x�z�p�Z��T�ƅ�@��C�����x�x�x�x�z�p�Z��T�����r+��6���e�4�
�1�!�h����
����l������;�u�c�����������Z��h �����f�_�u�u�8�)����Q���F������u�u�u�u�w�}�W��Y����l�N��Uʴ�9�0�u�u�w�}�W���Y�����\�����u�u�u�
�/�.��������F�S����4�<�y�u�w�}�Wϭ�����R9��V��U���u�h�u�
�3�)�[���Y�����O�����4�<�u�u�w�`�W�������l�N��Uʦ�4�<�
�
�3�)�W���Y�����S��Y���u�u�u�8�6�4�(�������E��SN��U���#�9�1�_�w�}�W���&����l��B�����4�u�k�'�#�<����Y����9F�C�X���x�x�x�x�z�p�Z���
����^��C�X���x�x�x�x�z�p�Z���YӇ��XF�N�U���n�u�u�4�;�8�W���DӅ��9F������1�i�u�d�l�}�WϿ�����F�F��ڊ���x�u�8�3���D���O��_��]±�;�
� �d�j�u����&����{K��S�����u�k�r�r�~�}�����֓�F ��
N�����
���x�w�2����I���3�G�����1�;�
� �f�W�W���&����Z�
N��R�ߊu�u�
�1�#�}�K�������d/��C����!�u�u�k�p�z�W�������Z��U��U���u�<�d����FϺ�����F�I��\���:�u�1�;��(�F��Qӂ��9��s:��Dʱ�"�!�u�u�i�z�P���Y������1����u�u�1� �w�}�W������G��=N��U���x�x�x�x�z�p�Z��T�ƅ�C��U�����x�x�x�x�z�p�Z��T�����T��U¶�>�u�0�<�]�}�W���Y����_��A��U���u�9�u�u�f�}����Y���F�N��ʶ�u�u�d�u�?�3�W���Y���F�N�����7�3�u�h�3�3�L���Y���F�N��U���d�7�3�u�j�9���Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�0�1�6�>��������9