-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���lǶd�����,�<�0�n�]�.�W���ݕ��l
��^��D��4�9�u� �2�4��������T��B �����{�9�n�_�9�4�ϳ�<����p ��1�����d�a�
�4�w�.�}���Y����A��=N��U���u�u�u�0��$����Y�ƿ�A��T��W���6�w�u�u�w�}�W���Yӂ��W��N��Oʼ�!�2�'�o�w�o�W���Y���F������u�u�o�<�#�:���Y���F�N��U���8�8�&�/�w�}�MϷ�����\�d��U���u�u�u�%�%�}�}���Y���F��S�U���o�<�u�!��2����������S��Dʱ�"�!�u�|�w�}�W���Y����VV�N��U���;�&�1�9�0�>�W���Y���F��N��U���u�u� �u�#�����&����\��@����1�"�!�u�~�W�W���Y���R��N��U��<�u�!�
�8�4�(�������D��_C����!�u�|�u�w�}�W���YӅ��F�N��U���&�1�9�2�4�}�W���Y�����N��U���u�;�&�1�;�:��������W��C��U���;�:�e�n�]�}�W���Y�ƻ�F�N��Oʼ�u�!�
�:�>�f�}���Y���F��N��U���o�:�!�&�3�1��������AN��^
��X���:�;�:�e�l�}�W���Y����_�N��U��<�u�!�
�8�4�W���Y����9�������u�_�4�6�>�8����Y����\ ��+��Dۖ�3�e�7�3�g�l�Cց��ƥ�l��^	��ʴ�1�e�!�%�m�.��������V��EF�����x�u�:�;�8�m�L���������E_�����u�!�
�:�>�����ۇ��W��N�����u�|�u�!�'�}��������Z��E��U��!�u�0�
�>�8�F���ӕ��l
��^�����'�}�"�1�?�l��������F��_��ʣ�'�4�9�u�6�}�W���&����J]ǑV�����0�&�;�'�:�)����Y����]��=�����!�u�,�
�6�.�����ƾ�^F��A�����u�&�w�9�4�����s����Z��RN�����,�0�o�&�%�3�L������G��V�����u�3�'�8�m�+�����ƥ���h�����!�'�7�!�w��>���<����v!��c+��'�����o�&�%�3�L�������9l��R�����6�&�
� �%��MϮ�����N��S�U��2�;�u�u�w�<�������F��S����,�!�0�<�w�/��������Ul�N�������
����_��������h����u�=�;�u�w�}�W���Y����9��GN�Uº�=�'�u�k�p�z�L���Y����_��=N��U���u�u�4�1�g�)���Y����]ǻN��U���u�3�_�x�.�)����Y����@
��R1�����u�'�6�&�l�W�(�������P��D1�U���6�&�u�6�<�}�}�����ƹF��QN�����#�;�u�;�w�1�W���H����[��N��U���<�u�6�e�j�z�P������F�N��U���$�u�h�'�:��9���7����aN��S�����|�u�u�u�w�}������ƹF��Y
�����;�u�'�6�$�f�}�������P��D1�����d�u�'�6�$�}����H����V��=N��U���1�'�
�8�w�`����H���@��_��ʡ�4�&�4�0�8�;�W���Yӏ��%��a1��!����4�1�d�w�}�������F��R ךU���u�u�u�4�3�l����E����G��DN��U��|�_�u�u�w�1��ԜY���F���ۊ�8�u�h�4�3�l�}���Y�Ʃ�WF��d����=�&�&�!�6�.�������WF��X���ߠ%�8�8�'��>����H�Ƽ�\��DN�����u�7�2�;�]�}�W���Q����V��CN��ʶ�>�h�r�r�w�5����Y�������U���d�|�!�0�w�}�W���Y�������U���d�|�!�0�w�}�W���Y���F���]��������<�������\�S_����u�u�u�u�w�3�W���s���F�N�����h�'�8����9���<�έ�W��C��\���u�u�u�u�2�9���Y����]��QU�����'�6�&�n�]�8�Ϭ���Ɠ��V��<���n� �0���s��������W����N���;�<�,�8���F���&ù��U9��\�U���u�u�2�;�%�>�_���Y���"��V9�����u����w�`�D��Y���F��S
�����;�0�o����%��Y��ƹF�N�����&��1�=�m��#���+���O��N�����u�_�u�u�w�}����Y�ƅ�5��h"��<��u�u�u�u�4�6�Mϗ�Y����)��tUךU���u�u�1�'�$�m�Mϗ�Y����)��t1��6���}�1�'�&� �9���HӢ��}2��G�U���u�u�6�e�m��W���&����p]ǻN��U���e�o�����;���:����g)��s��"���=�x�d�� �	�W���s���F�V
�����u�u�����0���/����aN��S�����!�u�u�u���8��B���F���U���������}���Y���D��N��U���
���n�w�}�W�������z(��c*��:���
�����)� ������"��y:��E��u�u�u�u�&�}�W���Y����)��t1��6���}�4�4�<�#�}�W���6����V�d��ʰ�!�!�n�_�%�5��������A��X��C���d��3�e�5�;�G��M�ƥ�9F������;�u�c��f���������lW��1��ʼ�_�u�u�u�w�2����Y���F�N�����u������4�ԜY���F�N����o��u����>���<����l�N��U���u�6�e�o��}�#���6����9F�N��U���u�e�o����3���>����v%��eUךU���u�u�u�u�3�/�W���7ӵ��l*��~-��0����_�u�u�w�}�W�������z(��c*��:���n�u�u�u�w�}�WϺ�Y�ƅ�5��h"��<������_�w�}�W���Y�ƻ�F��~ ��!�����n�u�w�}�W���Yӗ��	F��cN��1��������t�}���Y����P	��X ���ߠ_�7�2�;�w�}�ٛ�;�׏�U9��U��E��a�
�4�
�w�}����������u,�6���e�7�3�e�f�i�(���s���C	����U�ߊu�u�u�u�;�}�IϽ����F�N����h�u�1�'�$�m�}���Y���P��
P�����u�u�u�u�&�}�Iϯ�U���F������k�4�1�0�$�q�W���Y����VW�	N��D�ߊu�u�u�u�f�`�W��s���F�@�H���0�y�u�u�w�}����Gӗ��l��Y
�����!�6� �0�]�W