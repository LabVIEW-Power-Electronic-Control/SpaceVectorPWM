-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ��m�d�a���(���
����GF�N�����9�u�u����;���:���F��h��U���������}���Y����G��T��;ʆ�����]�}�W�������	F��cN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�%�<���6����g"��x)��N���u�<�
�9�?��W���7ӵ��l*��~-��0����}�d�1� �)�W���s���Z��V��U���������!���6���F��@ ��U���_�u�u�;�5�)�(���Y����g"��x)��*�����}�d�3�*����P���F��h�� ���e�o�����;���:����g)��]����!�u�|�_�w�}��������F��x;��&���������W��Y����G	�UךU���%�'�!�'��}�W���Y����)��t1��6���u�f�u�:�9�2�G��Y����C9��T��;ʆ�����~�W���s����[��T��ʷ�=�#�:�u�e�e�Fޚ��֓�lW��DNךU���:�&�4�!�6�����&����P9��N��1�����o�u�f�f�W�������R��V�����
�:�<�
�w�}�#���6����	[�I�U���6�;�!�;�w�-�$���¹��^9��N��1��������}�E�������V�S��E��e�e�e�e�g�m�G��H��ƹF��X �����4�
��&�e�;���Cӵ��l*��~-��0����}�e�1� �)�W���C���V��^�E��e�e�e�d�u�W�W�������]��G1��*���
�&�
�u�w�	�(���0����p2��F�U���;�:�e�u�j��G��I����V��^�D��n�u�u�6�9�)����	����@��Q��F��������4���Y����W	��C��\��u�e�e�e�g�m�G��I����V�=N��U���&�4�!�4��	��������\��c*��:���
�����m��������\�^�E��e�e�e�e�g�m�G���s���P	��C��U����
�!�
�$��W���-����t/��a+��:���g�u�:�;�8�m�W��[����V��^�E��e�e�e�n�w�}��������R��c1��B���8�c�o����0���/����aF�N�����u�|�o�u�g�m�G��I����W��^�W�ߊu�u�:�&�6�)����-����l ��hY��U���
���
��	�%���Iӂ��]��G��H���e�e�e�e�g�m�F��I����l�N�����;�u�%���)�(���&����`2��{!��6�����u�g�w�2����I����D��^�E��e�d�e�e�g�m�L���YӅ��@��CN��*���&�d�
�&��}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��_�E��e�e�n�u�w�>�����ƭ�l5��D�*���
�e�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�W�ߊu�u�:�&�6�)����-����9��Z1�U����
�����#���Q����\��XN�U��w�e�e�e�g�l�G��I����D��N�����!�;�u�%����������F��d:��9�������w�o�W������F��L�E��e�d�e�e�g�m�G��B�����D��ʴ�
��&�d��.�(��Cӵ��l*��~-��0����}�e�1� �)�W���C���V��^�E��e�e�e�e�u�W�W�������]��G1��*���`�3�8�d�w�}�#���6����e#��x<��G���:�;�:�e�w�`�U��I����V��^�E��e�n�u�u�4�3����Y����g9��X�����`�o�����4���:����T��S�����|�o�u�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
����U��X��U���
���
��	�%���Iӂ��]��G��H���e�e�e�e�g�m�G��I����l�N�����;�u�%���)�O�������	F��s1��2������u�e�}�������	[�^�E��e�e�e�e�g�m�G��Y����\��V ������&�d�
�$��O��*����|!��h8��!���}�e�1�"�#�}�^��Y����V��^�E��e�e�e�w�]�}�W���
������d:�����3�8�d�u�w�	�(���0����p2��F�U���;�:�e�u�j��F��I����V��^�E��n�u�u�6�9�)����	����@��h��*��o������!���6���F��@ ��U���o�u�d�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lV�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
����9��N��1��������}�GϺ�����O�
N��W�ߊu�u�:�&�6�)��������_��h[��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�E���_�u�u�:�$�<�Ͽ�&����G9��\��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�D��w�_�u�u�8�.��������]��[�*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��d�d�w�_�w�}��������C9��Y����
�g�o����0���/����aF�N�����u�|�o�u�g�m�G��I����V��^�E��e�d�e�e�l�}�WϽ�����GF��h�����#�g�d�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�f�f�W�������R��V�����
�#�g�g�m��3���>����v%��eN��Dʱ�"�!�u�|�m�}�G��I����V��^�E��e�e�e�e�g�m�L���YӅ��@��CN��*���&�
�#�g�a�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�l�G��Y����\��V �����:�&�
�#�e��Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�m�F��B�����D��ʴ�
�:�&�
�!�o�F���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��H����F�T�����u�%�6�;�#�1�D݁�Y�Ɵ�w9��p'��#����u�f�u�8�3���Y���V��^�E��e�e�e�e�g�m�G��I����l�N�����;�u�%�6�9�)���&����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������V�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����W��^�����u�:�&�4�#�<�(���
���� T��q_��0��o������!���6���F��@ ��U���o�u�e�d�f�l�G��I����V��_�E��e�e�n�u�w�>�����ƭ�l��D�����f�m�e�e�w�}�#���6����e#��x<��F���:�;�:�e�w�`�U��H����V��^�E��e�e�e�e�g�m�U�ԜY�Ư�]��Y�����;�!�9�f��i�Mύ�=����z%��r-��'���d�1�"�!�w�t�M���I����V��^�E��e�e�e�e�g�l�F��B�����D��ʴ�
�:�&�
�!�o�F���Y����)��t1��6���u�f�u�:�9�2�G���D����V��^�E��e�e�e�e�g�m�G��H����F�T�����u�%�6�;�#�1�D݁�<����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��H����]ǻN�����4�!�4�
�8�.�(���&���5��h"��<������}�w�2����I����D��_�D���_�u�u�:�$�<�Ͽ�&����G9��]��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������V��^�U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�E��w�_�u�u�8�.��������]��[��E��������4���Y����\��XN�U��w�e�n�u�w�>�����ƭ�l��D��ي�u�u��
���(���-���F��@ ��U���o�u�d�d�l�}�WϽ�����GF��h�����#�
�u�u���8���&����|4�N�����u�|�o�u�f�m�L���YӅ��@��CN��*���&�
�#�
�w�}�#���6����e#��x<��Gʱ�"�!�u�|�m�}�F��B�����D��ʴ�
�:�&�
�!��W���-����t/��a+��:���g�1�"�!�w�t�M���H���9F������!�4�
�:�$��ׁ�Y�Ɵ�w9��p'��#����u�b�1� �)�W���C���V��^�N���u�6�;�!�9�}��������EW��^�U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��[���F��Y�����%�6�;�!�;�l�(��I����g"��x)��*�����}�a�3�*����P���W��_�E��e�e�w�_�w�}��������C9��Y����
�e�u�u���8���&����|4�Z�����:�e�u�h�u�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������V��N��1��������}�F�������V�S��E��e�d�e�e�g�m�L���YӅ��@��CN��*���&�
�#�`�c�m�Mύ�=����z%��r-��'���a�1�"�!�w�t�M���I����V��^�E���_�u�u�:�$�<�Ͽ�&����G9��X��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�����u�:�&�4�#�<�(���
���� R��q(��3���u�u��
���(���-��� U��X����u�h�w�d�f�l�F��H����W��_�D��d�d�d�w�]�}�W���
������T�����f�
��o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�d�d�f�m�L���YӅ��@��CN��*���&�
�#�a�f�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��B�����D��ʴ�
�:�&�
�!�o�@���I����	F��s1��2������u�d�}�������	[�_�D��d�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������F��d:��9�������w�n�W������F��L�E��e�e�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-��������lT�=��*����
����u�W������F��L�E��n�u�u�6�9�)����	����@��A[��U����
�����#���Q�ƨ�D��^��O���e�e�d�n�w�}��������R��X ��*���
�u�u����>���<����N��S�����|�o�u�e�f�m�L���YӅ��@��CN��*���&�
�#�
�w�}�#���6����e#��x<��Eʱ�"�!�u�|�m�}�G��s���@��V�����
�&�u�u���8���&����|4�^�����:�e�u�h�u�m�G��I����V��^�D��u�u�4�!�>�(�ϸ�����\��PN����;�n�u�u�6�)����Ӏ��l��X
��ʺ�u�%��
�$�}�W�������@F��X ��N���u�&�2�4�w�-��������`2��C_�����u�u��
���L���Yӕ��]��V�����1�
�l�o���2���s���@��V����� �l�
�g�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������V��]��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�'�.��������l��h��*���u��
���f�W���
����_F��h��*���
�e�o����9�ԜY�ƿ�T�������6�0�
��$�l�(���&���5��h"��<��u�u�&�2�6�}��������lP��N��:����_�u�u�>�3�Ϭ�����\��c*��:���
�����l��������l�N�����u�%�&�2�4�8�(���
�ߓ�@��T��!�����n�u�w�.����Y����Z��S
��L������]�}�W�������C9��P1������&�d�
�$��F��*����|!��d��Uʦ�2�4�u�%�$�:����A����q)��r/�����u�<�;�9�6�����
����g9��W�����m�o�����4�ԜY�ƿ�T�������7�1�l�u�w��;���B�����Y������-� �
�b����K����	F��s1��2������u�d�}�������9F������3�
��-�"��Bځ�����Q�=��*����
����u�FϺ�����O��N�����4�u�%�&�0�>����-����l ��h_��U���
���n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��h�����
�:�<�!�1��Bہ�H����g"��x)��*�����}�d�3�*����P���F��P ��U���4�%�4�d�#���������T�=��*����
����u�FϺ�����O��N�����4�u�8�
��(�F���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�
�0�
�e�j�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������A��\�U����
�����#���Q�ƨ�D��^����u�<�;�9�1��5�������9��C����� �d�e�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����U5��u=�� ���`�
�
�:�>�)����H����	F��s1��2������u�d�}�������9F������!�%�d�
�"�o�N���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����a�'�2�d�g�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h��D���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����A��]�U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-����&����CT�=��*����
����u�W������]ǻN�����9�!�%�&�%�:�F��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����2�6�0�
��.�D������5��h"��<��u�u�&�2�6�}��������lW��T��:����n�u�u�$�:����*����
^��h��@���%�u�u����>���<����N��
�����e�n�u�u�$�:����*����
^��h��*��d�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�&����_��h��@���%�u�u����>���<����N��
�����e�n�u�u�$�:����*����W��1����g�u�u����>���<����N��
�����e�n�u�u�$�:����*����W��1��*��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������lW��hZ�����f�d�o����0���/����aF�N�����u�|�_�u�w�4��������lW��hZ�� ��a�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G9��1�����d�f�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����\��h��C���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϱ�&����9��P1�A���u��
����2���+����W	��C��\�ߊu�u�<�;�;�.����	�ӓ�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�$�1����L����lW��N�&���������W������\F��d��Uʦ�2�4�u�0��0�F؁�����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�l�(���&����\��c*��:���
�����}�������9F������&�9�!�%�n�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʦ�9�!�%�l�%�:�F��Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V����� �l�
�g�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������`9��s*�� ���c�
�0�
�d�d�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��G1�����0�
��&�`�;���Cӵ��l*��~-�U���&�2�4�u�'�.��������\��x!��4��u�u�&�2�6�}�$���,����|��X��F���
�m�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������`9��b"�����
�c�
�
�2��D��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����2�6�0�
��.�F܁�
����\��c*��:���n�u�u�&�0�<�W���
����W�� ]��U�����n�u�w�.����Y����G9��D�����!�'�
�d�n�;�(��&���5��h"��<������}�f�9� ���Y����F�D������6�
�4�2���������9��E��D��u�u��
���(���-��� W��X����n�u�u�&�0�<�W���
����@��d:�����3�8�d�u�w�	�(���0��ƹF��^	��ʴ�
�<�
�1��e�W���6����}]ǻN�����9�3�
�!��.�(�������V9��hW�� ��m�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G9��D�����!�'�
�m�n�/���@����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�
�!��&��)��������l^��B1�@���u�u��
���(���-��� W��X����n�u�u�&�0�<�W�������@��C�����
�`�m�'�0�l�G���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N����
�0�:�2�9�;�(��J����	F��s1��2������u�g�9� ���Y����F�D�����8�
�b�1�:�/��������^�=��*����
����u�W������]ǻN�����9�!�%�f��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʡ�%�f�
�0��i�D��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��D�����c�
�0�:�0�3����I�ޓ�F��d:��9�������w�m��������l�N�����u�0�
�8�f�k��������A��Z�U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�Eځ�����R��B1�Mފ�g�o�����4���:����V��X����n�u�u�&�0�<�W���&�ӓ�V��P�����d�g�u�u���8���&����|4�N�����u�|�_�u�w�4��������9��h_�G���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����J˹��T9��V��U���
���
��	�%���Y����G	�UךU���<�;�9�&�;�)���&����A��h��D��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CW��h
�����;�'�2�d�d�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h]�����'�4�
� �f�i�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
�0�:�2�9�/���J����`2��{!��6�����u�e�3�*����P���F��P ��U���
�f�3�
�f�n����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���'�2�d�a�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�C���8�'�4�
�"�l�@߁�K����g"��x)��*�����}�u�8�3���B�����Y�����!�%�m�
�2�2��������R��N��1��������}�GϺ�����O��N�����4�u�'�
�"�d�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V����� �l�
�d�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������C9��P1������&�a�3�:�n�Mύ�=����z%��N�����4�u�%�&�0�?���O����|)��v �U���&�2�4�u�'�.��������l��1����o������}���Y����R
��G1�����1�g�f�o���2���s���@��V�����2�6�0�
��.�Fہ�
����\��c*��:���n�u�u�&�0�<�W���
����W��^��U�����n�u�w�.����Y����Z��D��&���!�b�3�8�f�}�W���&����p]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�2�'�;�(���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʲ�%�3�
�b�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h/�����
�`�
� �f�o����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*���-� �
�`��(�F���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʲ�%�3�
�e��m�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��E�� ��m�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����Z��D��&���!�d�3�8�e�}�W���&����p]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�2�'�;�(��&���5��h"��<������}�f�9� ���Y����F�D�����'�
� �d�c�-�W���-����t/��a+��:���f�u�:�;�8�m�L���Yӕ��]��P�����d�
�e�o���;���:����g)��]����!�u�|�_�w�}����Ӏ��r$��x�����
�a�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������A��B1�L���u�u��
���(���-��� W��X����n�u�u�&�0�<�W���8����F��[��*���g�l�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��h_�*��o������!���6�����Y��E��u�u�&�2�6�}��������l��N��1��������}�GϺ�����O��N�����4�u�'�
�"�l�O���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V����� �d�l�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������^��B1�M���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����H����P��G_��U���
���
��	�%���Kӂ��]��G�U���&�2�4�u�8�/����&����CT�=��*����
����u�W������]ǻN�����9�;�!�=��(�F���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�e�3�
�n��C��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��Dي� �g�f�%�w�}�#���6����e#��x<��G���:�;�:�e�l�}�Wϭ�����]	��_�����d�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����[��Q��E݊�g�o�����4���:����V��X����n�u�u�&�0�<�W���8����F��]����� �g�a�%�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����G�� 1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:����*����K)��h_�*���g�l�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�l'��O!��*���
�0�
� �e�m����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N����
� �g�c�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W������� ��v,��:���d�`�g�3��k�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V��&�����!�!��3�(���K�ѓ�F��d:��9�������w�n�W������]ǻN�����9�3�
��/�(�(݁�����l ��W�����u��
����2���+������Y��E��u�u�&�2�6�}����@����^��GZ��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�o�(���K�ד�F��d:��9�������w�o�W������]ǻN�����9�;�!�=�c�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʻ�!�=�a�3��l�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N����
� �g�l�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h\�����e�
�d�o���;���:����g)��\����!�u�|�_�w�}����ӈ��A��h��F���%�u�u����>���<����N��S�����|�_�u�u�>�3�ϰ�����l ��]�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����S��N�&���������W������\F��d��Uʦ�2�4�u�8��i����M����\��c*��:���
�����}�������9F������!�%�g�
�"�n�N���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����-���!�f�m����Lƹ��\��c*��:���
�����}�������9F������7�:�
��g�(�(��&����W��N�&���������W������\F��d��Uʦ�2�4�u�:�;�%�2ߑ�����l ��\�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)���&����W��N�&���������W������\F��d��Uʦ�2�4�u�8��l����O¹��\��c*��:���
�����}�������9F������<�8�
� �d�d����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���f�`�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:��������CT��B1�F���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������9��hZ�*��o������!���6���F��@ ��U���_�u�u�<�9�1����&����U��]��G��������4���Y����\��XN�N���u�&�2�4�w�0�(ׁ�����l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�k����Mʹ��\��c*��:���
�����}�������9F������&�9�!�%��(�C���	����`2��{!��6�����u�e�3�*����P���F��P ��U���6�
�m�g�1��Eց�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�8�c�1�:�/��������l��N��1��������}�GϺ�����O��N�����4�u�0�
�:�l�(�������l ��X�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�)��������9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-����Nǹ��\��c*��:���
�����}�������9F������&�9�!�%��(�C���	����`2��{!��6�����u�e�3�*����P���F��P ��U���6�
�m�f�1��Aށ�J����g"��x)��*�����}�d�3�*����P���F��P ��U���
�8�g�
�2�2�������� 9��T��!�����
����_�������V�=N��U���;�9�&�9�#�-�(���M�ߓ�F��d:��9�������w�m��������l�N�����u�0�
�8�o�;�(��&���5��h"��<������}�w�2����I��ƹF��^	��ʳ�
�!�l�
��(�C���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�
�!�d�l�1��Fׁ�J����g"��x)��*�����}�d�3�*����P���F��P ��U���6�
�d�
��(�B���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�
�!�d�l�d�;�(��&���5��h"��<������}�f�9� ���Y����F�D������6�
�d��(�B���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʳ�
�!�d�g�e�;�(��&���5��h"��<������}�f�9� ���Y����F�D������6�
�d�����H����	F��s1��2������u�d�}�������9F������3�
�!�d�e�h����Oʹ��\��c*��:���
�����l��������l�N�����u��6�
�f��(���L�ғ� F��d:��9�������w�n�W������]ǻN�����9�3�
�!�f�d�@���&����CU�=��*����
����u�FϺ�����O��N�����4�u��6��l�(ׁ�����l��N��1��������}�D�������V�=N��U���;�9�3�
�#�l�N�������9��T��!�����
����_������\F��d��Uʦ�2�4�u�8��o����K¹��\��c*��:���
�����}�������9F������<�8�b�3��o�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����;�!�3�
�c��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��C��D؊� �c�d�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������V
��Z�*���c�f�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��_�����'�4�
� �a�h����Y����)��t1��6���u�e�1�"�#�}�^�ԜY�ƿ�T����*���d�
� �c�f�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R����f�1�8�'�6����J����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�d��(�A���	����`2��{!��6�����u�e�3�*����P���F��P ��U���-��,� ��9�(��&����W��N�&���������W��Y����G	�UךU���<�;�9�9�4�����Iƹ��\��c*��:���
�����}�������9F������9�6��d�1��Fځ�H����g"��x)��*�����}�g�3�*����P���F��P ��U���
�
�
�f�1��Eځ�K����g"��x)��*�����}�u�8�3���B�����Y�����<�<�3�
�f��E��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��E�����3�
�f�
�d�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������hY�����3�
�f�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����@��C��*���b�d�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����ӕ��l��^�� ��b�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������l��h�����&�
� �b�b�-�W���-����t/��a+��:���d�u�:�;�8�m�L���Yӕ��]��D�����
� �b�f�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��e�����
� �b�d�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h��9����!�d�d�>�����&¹��lQ��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�#�-�D���&����CT�=��*����
����u�W������]ǻN�����9�!�%�`�1��Gށ�K����g"��x)��*�����}�u�8�3���B�����Y�����g�
� �m�`�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��Z��L���
�g�
�f�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƹ�C9��h��M���%�u�u����>���<����N��S�����|�_�u�u�>�3�Ϫ�	����U��]��F��������4���Y����\��XN�N���u�&�2�4�w��F���H����W��G]��U���
���
��	�%���Kӂ��]��G�U���&�2�4�u�:��@���&����CU�=��*����
����u�GϺ�����O��N�����4�u�
�0�"�)�Fށ�����l��N��1��������}�D�������V�=N��U���;�9�3�
���E�������l��Q����� �b�f�%�w�}�#���6����e#��x<��D���:�;�:�e�l�}�Wϭ�����@��C��D���
�c�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����ƿ�_9��G_�����b�
�g�o���;���:����g)��^�����:�e�n�u�w�.����Y����G��1��*��
�g�o����0���/����aF�
�����e�n�u�u�$�:����*����2��x��D���3�
�c�
�f�g�$���5����l0��c!��]��1�"�!�u�~�W�W������� ��T������'�6� �2�i�(݁�����l��N��1��������}�D�������V�=N��U���;�9�3�
�#���������F��_�� ��e�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����G9��D�����!�'�
�d�c�;�(��&���5��h"��<������}�f�9� ���Y����F�D������6�
�4�2���������9��Q��Gي�f�o�����4���:����U��S�����|�_�u�u�>�3�ϸ�&����R��d�����0�a�
� �o�j����Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*����&�
�!�"�)����A�ד�F9��1��U����
�����#���Q����\��XN�N���u�&�2�4�w���������G��C��*���g�3�
�a��n�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��d1��*���0��'�6�"�8�Cׁ�&����W��N�&���������W��Y����G	�UךU���<�;�9�3��)�4���&����P��R1�*���l�a�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�l��t��*��� �!�'�
�b�l����Oƹ��\��c*��:���
�����l��������l�N�����u��6�
�6�8�$�������lS��1��*��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������l%��R1����� �0�`�
��(�N���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʥ��9�
�
�"�d�D���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y������g�3�
�n��C��*����|!��h8��!���}�u�:�;�8�m�L���Yӕ��]��[��#���3�
�e�b�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��G1��ۊ� �d�d�
�e�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��^1��*���3�
�e�b�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������E��*���d�f�
�g�m��3���>����v%��eN��U���;�:�e�n�w�}�����Ƣ�G
��1��*��l�%�u�u���8���&����|4�N�����u�|�_�u�w�4��������F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�'��݁�&����S��G_��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�8��(ہ�����9��T��!�����
����_�������V�=N��U���;�9�9�6��h����I�ޓ�F��d:��9�������w�o�W������]ǻN�����9�!�%�<�>����N����\��c*��:���
�����}�������9F������!�%�<�<��h����I�ޓ�F��d:��9�������w�m��������l�N�����u�:�'�&��(�F��&���5��h"��<������}�w�2����I��ƹF��^	��ʻ�!�=�m�3��m�G���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V����� �d�f�%�w�}�#���6����e#��x<��Eʱ�"�!�u�|�]�}�W�������l0��1�����d�`�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ơ�P9��1��*��l�%�u�u���8���&����|4� N�����u�|�_�u�w�4��������lQ��B1�Gӊ�d�o�����4���:����T��S�����|�_�u�u�>�3�Ϫ�	����9��h_�F���u�u��
���(���-���F��@ ��U���_�u�u�<�9�1��������P��B1�Fӊ�g�o�����4���:����V��X����n�u�u�&�0�<�W�������U��[�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�3����H����W��h�Oʆ�������8���Iӂ��]��G�U���&�2�4�u�%����A����	F��s1��2������u�g�9� ���Y����F�D�����0�
�8�g��(�F��&���5��h"��<������}�f�9� ���Y����F�D������!�'�d������&����p	��T��*���d�b�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������V
��Z�*���d�e�
�f�m��3���>����v%��eN��Dʱ�"�!�u�|�]�}�W�������`9��E��<���4�2�
�;��2����O����W��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�$�1����K����T��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�1�����&����R��h��*���'�0�c�d�1��E���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʺ�!� �0�6�9��(�������@��h��D��
�f�o����0���/����aF�N�����u�|�_�u�w�4��������C��R ��A���<�0�4�&�0����H¹��\��c*��:���
�����l��������l�N�����u� �
�%�%�8��������l��^	�����d�e�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƫ�C9��hW�����u��
���f�W���
����_F��h��*���$��
�!��.�(���Y����)��tUךU���<�;�9�4��4�(���&����	F��x"��;�ߊu�u�<�;�;�:����&�ѓ�VF��d:��9����_�u�u�>�3�Ϲ�	����V��X�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�:����&����\��S��U���
���
��	�%���Y����G	�UךU���<�;�9�2�'�;�(��&����W�=��*����
����u�W������]ǻN�����9�4�
��1�0�Mύ�=����z%��r-��'���e�1�"�!�w�t�}���YӅ��C	��Y��G��d��3�e�1�9�(���
����@9��h]�� ���1�%��_�w�}�������F�N��<���u����l�}�W���YӨ��l5��p+��U�����n�u�w�}�WϺ�ù��w2��N��!����_�u�u�w�}����.����\��y:��0��u�u�u�u�3�(�(���-����z(��p+��\�ߊu�u�:�!��}�W���YӅ��\��yN��1�����_�u�w�}�W�������z(��c*��:���n�u�u�u�w�9����Y����g"��x)��*�����}�d�3�*����P���F�N�����u������4���:����U��S�����|�_�u�u�w�}���0�Ɵ�w9��p'�����u�u�u�:�#�g�8���*����|!��h8��!���}�d�1�"�#�}�^���s���V��T�����!�_�_�u�w�2�����ơ�w^��*��*ڊ�8�9�f�;��o���&¹��K9��GN�����u�0�0�<�w�W�W���Y�ƅ�\��y:��0��u�u�u�u���$���<����}2��r<�U���u�u�1�;���#���Y����t#��=N��U���u�<�d����Mϗ�-����l�N��Uʱ� �
���w�}�9���<���9F������u�u�u�u�3�3�W���7ӵ��l*��~-��0����}�d�1� �)�W���s���F�S��U���������!���6���F��@ ��U���_�u�u�u�w�2���6����g"��x)��*�����}�d�3�*����P����F�R �����:�0�!�_�]�}�W���	����GF��sV�D���
�
�6�%�d�3�(���
�ד�/��N�����'�6�}�u�w�}�Wϗ�Y�ƅ�g#��eUךU���u�u� �
���W���7����a]ǻN��U���<�e����g�>���>����F�N�����
���u�w��2���B���F�
�������o����%���s���C	��FךU���u�u�<�e�m��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����Z��N��U���
���
��	�%���Hӂ��]��G�U���u�u�:�6�3�}�W���*����|!��h8��!���}�u�:�;�8�m�L���Y�����CN�:���������4���Y����\��XN�U��u�u�0�1�4�0������Ɠ9��^ ךU���
�
�4�1�d�3�(���
���� 9��[�����e�o�6�8�8�8�ϳ�=����wR��1�����g�&�f�;��o�D�������Cl�N�����6�8�%�}�w�}�W���0���W�N��U��������`�W��Y���F��^ ��"����h�u�g�]�}�W���Y����l1��c&��K��y�u�u�u�w�9����0����X�GךU���:�!�8�%��}�W���YӅ��[�V�����u�u�u�u�%�.���Y����@�N��U���1�;�u�k�0�-����J����9F�N��U���d�h�u�'��(�N܁�H���F�N��U��2�%�3�
�d�>�[���Y�����CN��U���
� �l�
�e�f�}���Y����U��h]����;�
�g�f�1�1�(���&�����G�����g�m�d��1�m����&�Ԣ�lU��D1�*ي� �9�1�%�w�}��������R�=N��U���u��h�u�{�}�W���YӨ��l5��p+��K��_�u�u�u�w�4�G���=���F��d��U���u�1�;�
��	�W���J��ƹF�N��������h�w�o�}���Y������FךU���u�u�9�u�i�<�(���U���F������k�4�
�&�{�}�W���Yӂ��F�	��*���l�
�e�_�w�}�W������F��G1��*���%�y�u�u�w�}����GӁ��l ��Y���ߊu�u�u�u�8�)�J�������l_��G\����u�3�e�3�"��E���J���� T��h��*���
�g�o�6�:�2��������W��Q1�����
�g�&�f�9��E�������@ǻN�����<�u�4�u�]�}�W���Y���F��=N��U���u� �
���}�I��s���F�S��*����u�k�f�{�}�W���Yӂ��9��s:��H���g�_�u�u�w�}����.����[�\��U���%�'�u�4�w�W�W���Y�ƨ�]V�	N��*���-� �
�`��(�F���	��ƹF�N����h�u�������L����V��G_�U���u�u�1� �w�c����;����G9��1��*��
�g�n�_�w�}�(߁�������\��*ۊ�
�f�o�6�:�2��������W��Q1�����
�g�&�f�9��(�ԜY�ƫ�]��TN�����u�u�u�u��}�I��s���F�y;��&����h�u�y�w�}�W�������d/��N��U��_�u�u�u�w�4�F���=���F��d��U���u�1� �
��	�W���H���F��E�����_�u�u�u�w�4�G��Y����U��V��E�ߊu�u�u�u�>�l�J�������lW��h����u�u�u�%�8�8�J�������lW��h�����_�u�u�u�w�2���Y����U��V��G��_�u�u�
��>�������]��h_��A��6�8�:�0�#�0�3��H�Ҫ�9��Z��G���f�;�
�
�]�}�W�������^��d��U���u��u�k�f�W�W���Y�Ƃ�~9��v)��H���y�u�u�u�w�9�߁�0����X�BךU���u�u�<�d� ��?��Y����F�N�����
���u�i�l�}���Y������FךU���u�u�<�e�j�}��������l��=N��U���u�<�d�h�w�/�(���H�ғ�JǻN��U���%�:�0�h�w�/�(���H�ғ�C��RBךU���u�u�:�!�j�}��������l��dךU���
�
�6�%�d�3�(���
�ד�l3��N�����0�!�8��o�l�C���&����lU��D1����
�_�u�u�2�8�������F�N��<���k�d�_�u�w�}�W���&����vF�_�U���u�u�1�;���#���G����9F�N��U���d����j�}�E�ԜY���F��B��<���u�k�d�_�w�}�������9F�N��U���e�h�u�'��(�F���	��ƹF�N����h�u�'�
�"�l�N���U���F������h�u�'�
�"�l�N�������9F�N��U���!�h�u�'��(�F���	����9lǑ=N��U���!�0�6�'�2�)�����έ�l%��Q��U���!�0�&�4�2�0�������9F���6���&�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y����_��N��U���u�u�u�u�>�}�_�������l
��^��U���%�6�|�u�?�3�}���Y���F�N��U���4�
��3�:�a�W���7����^]ǻN��U���u�u�u�u�9�}����Y���F�N�����3�_�u�u�w�}�������F��SN�����&�_�_�u�w�p�����Ƽ�\��D@��X���u�%�:�0�$�u�������F��P��U���u�u�<�u�6���������R��V�����u�d�|�!�2�W�W���Y���F��F�����:�&�
�:�>��W���	������F��*���&�
�:�<��}�W���
����@��d:��؊�&�
�|�|�#�8�}���Y���F�N������-� �
�b��(�������V��W�I�������#�l�B�������G9��h_�*��_�u�u�u�w�}�W���Y����_��h_�����!�'�2�d�o�}�JϷ�&����R9��C����� �d�a�%�l�}�W���Y���F���*���'�2�d�e�w�`����Hǹ��lT��h����u�u�u�u�w�}�W���&�Г�V��^�I���'�
� �d�c�-�L���Y���F�N��U���
�
�0�
�e�j�K�������U��Z��G�ߊu�u�u�u�w�}�W�������A��\�U��2�%�3�
�g��E�ԜY���F�N��ʼ�n�u�u�u�w�8�Ϸ�B����������n�_�u�u�z�<����Y����V��C�U���%�:�0�&��-����s���Q��Yd��U���u�<�u�4��1�P����ƭ�WF��h��U���d�|�!�0�]�}�W���Y���Z �F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h_��U���6�|�4�1�9�)�_���
����[��G1�����9�2�6�e�~�t����s���F�N��U���3�
��-�"��Bځ�����Q�
N��*���-� �
�`��(�F���	��ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�w�}�Z���
������T��[���_�u�u�'�4�.�Wǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�r�r�w�5����Y���F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���f�3�8�g�~�}����Y���F�N��U����6�
�d������J���F��h��D���a�3�
�b��n�}���Y���F�N�����!�d�l�a�%�:�F��Y����`9��h_�*ފ� �c�a�%�l�}�W���Y���F������d�
�
�0��n�A��Y����G9��1�����f�
�f�_�w�}�W���Y���F��h��LҊ�
�0�
�f�f�a�W�������lR��B1�D���n�u�u�u�w�}�W���YӉ��P	��1����a�u�h�:��2�ށ�����l��=N��U���u�u�u�u�w�8�(���Hƹ��T9��V��Hʦ�9�!�%�`�1��Bց�K���F�N��U���u�&�9�!�'�j����H����[��R����
� �c�b�'�f�W���Y���F�N�����8�d�
�0��n�E��Y����G��1��*��
�g�_�u�w�}�W���Y���G��D1����d�u�h�!�'�.����I����l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�e�3�:�l�^�������F�N��U���u�u�3�
�#���������F��_��*���
�f�e�i�w���������G��C��*���l�3�
�f��n�}���Y���F�N�����!��&�
�#�(����&�ޓ�l��h_�C��u��6�
�6�8�$�������lR��1��*���
�f�_�u�w�}�W���Y���U5��C1�����!� �!�'��h�O�������F������4�0��'�4�(���&˹��l_��h����u�u�u�u�w�}�W���&����P��R�����'�2�d�d�w�`��������9��Z����� �d�a�
�e�W�W���Y���F�N�����%�b�
�0�8�:�������� F���*���d�c�1�8�%�<�(���H����CT��N��U���u�u�u�u�$�1����AŹ��^	��V �����a�m�i�u�2����O����\��Y1��*��e�%�n�u�w�}�W���Y�����h_�����'�4�
�0��i�O��Y����Q��R�����3�
�e�f�'�f�W���Y���F�N�����`�1�8�'�6�����M���F��G1�*���:�2�;�3��m�C���B���F�N��U���u�8�
�f�3�0����&����R��R�����f�
�0�:�0�3����H�ӓ�]ǻN��U���u�u�u�u�:��D������� F���*���3�
�e�d�'�f�W���Y���F�N�����m�'�2�d�e�}�JϪ�	����U��^����u�u�u�u�w�}�W������� 9��P1�A���h�!�%�a��(�F��&����F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W������]F��X�����x�u�u�%�8�8����	����l�N�����u�u�u�u�>�}��������V��V �����9�u�u�d�~�)��ԜY���F�N��U���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�t����s���F�N��U���3�
����)�F������� P��S����� �l�
�g�]�}�W���Y���V��^�U���u�u�0�1�>�f�W�������A	��D����u�x�4�&�0�}����
���l�N�����&�}�%�6�<�W�W�������F�N�����4�
�9�r�!�3�W���Y����_�I�\ʡ�0�_�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���|�!�0�_�w�}�W���Y���F��h��9����!�d�d�d�/���N��� ��O#��!ػ� �
�c�
��(�O���	��ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�w�}�Z���
������T��[���_�u�u�'�4�.�Wǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�r�r�w�5����Y���F���]���4�
�:�&��2����Y�ƭ�l����U´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�}��������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����Г�@��G��\ʡ�0�_�u�u�w�}�W���Y�ƾ�T9��N�U���
� �l�
�e�W�W���Y���F��SN��N���u�u�u�0�3�4�L���YӃ����T��N�ߊu�u�x�4�$�:�W�������K��N�����0�&�}�%�4�6�}���Y����]l�N��Uʼ�u�4�
�9�p�+�����ƭ�l��S��D���!�0�_�u�w�}�W���Y���N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��1����|�:�u�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�f�����H����AF�V�����
�:�<�
�w�}����PӇ��N��h�����:�<�
�u�w�-��������`2��C_�����d�|�|�u�?�3�W���Y���F�N�����a�u�h�2�'�;�(���	��ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�w�}�Z����Ƣ�K��C��U´�
��3�8�w�;����
������_��[���_�u�u�%������
����l��TN����0�&�}�%�$�<����	����U�������u�u�7�2�9�}�W���YӅ��VF��h-�����<�_�u�u�w�}�W�������C9��h��*���
�u�k�_�w�}�W���Y���F��F�����:�&�
�:�>��W���	������ ��]´�
�!�'�u�w�-��������Z��G��U���;�u�u�u�w�}�W���Y�����y=�����h�4�
��$�o����H���F�N��U���u�0�&�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�u�u�9�}��ԜY���F�N�����%��
�!��.�(���G���F�N��U���u�<�u�}�'�>��������lW������u�=�;�u�w�}�W���Y���F���;���&�u�h�4��	��������l�N��U���u�u�u�0�$�W�W���Y���F�N��Uʴ�
��3�8�k�}����&����U��UךU���u�u�u�u�w�}�������F�N��Uʢ�0�u�%���)�(���&���l�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U����
�&�u�j�<�(���
�ғ�@��d��U���u�u�u�u�w�8��ԜY���F�N��U���u�4�
��1�0�K���	����@��Q��G�ߊu�u�u�u�w�}�W����ƥ�l�N��U���u�"�0�u�'��(���&���� F�d��U���u�u�u�u�w�4�W���	����@��X	��*���u�%�6�|�w�5����Y���F�N��U���u�%��
�$�}�JϿ�&����GS��D��N���u�u�u�u�w�}�Wϻ�
���F�N��U���u�u�u�4������E�ƭ�l5��D�����f�_�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�"�2�}����&����U��N��U���u�u�u�u�w�}�WϷ�Y�έ�l��D�����
�u�u�%�4�t�W������F�N��U���u�u�u�%������DӇ��`2��CX�����n�u�u�u�w�}�W���YӃ��Vl�N��U���u�u�u�u�w�<�(������F��h=�����3�8�a�_�w�}�W���Y���F��SN��N���u�u�u�u�w�*����	����@��Q��@��u�u�u�u�w�}�W���Yӏ��N��h�����:�<�
�u�w�-����Y����9F�N��U���u�u�u�u�w�-�9���
�����d:��݊�&�
�n�u�w�}�W���Y�����Rd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�c�3�8�b�W�W���Y���F�N��ʼ�n�u�u�u�w�}�Wϩ��ƭ�l5��D�����c�h�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���7����^F���&���!�
�&�
�l�}�W���Y���F������u�u�u�u�w�}�W���YӇ��}5��D��Hʴ�
��&�b�1�0�A�ԜY���F�N��Uʰ�1�<�n�u�w�}�W���Yӑ��]F��h=�����3�8�b�h�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���0�u�u�u�w�}�W���Y�����y=�����h�4�
��$�e����N���F�N��U���u�0�1�<�l�}�W���Y�����YN��*���&�l�3�8�o�`�W���Y���F�N��U���}�4�
�:�$�����&���R��RG�����_�u�u�u�w�}�W���Y���R��d1����u�%��
�#�m����@���F�N��U���u�0�&�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�u�u�9�}��ԜY���F�N�����%��
�!�g�;���D��ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���H����lW��=N��U���u�u�u�u�w�1����Y���F�N��U���u�%��
�$�}�JϿ�&����GW��Q��L�ߊu�u�u�u�w�}�W����ƥ�l�N��U���u�"�0�u�'��(���H����lW��
P��U���u�u�u�u�w�}����Q����\��h�����u�u�%�6�~�}����Y���F�N��U���u�u�%���.�W������l��1����n�u�u�u�w�}�W���YӃ��Vl�N��U���u�u�u�u�w�<�(������F��h=����
�&�
�e�]�}�W���Y���F�R ����u�u�u�u�w�}� ���Y����g9��\�����d�h�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W������G��=N��U���u�u�u�u�w�}�W���7����^F���&���!�f�3�8�f�f�W���Y���F�N�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�f�����H���F�N��U���u�0�1�<�l�}�W���Y�����YN��*���&�d�
�&��o�J���Y���F�N��U���3�}�4�
�8�.�(�������F��h��\ʡ�0�_�u�u�w�}�W���Y���F��h �����i�u�%���)�C�������9F�N��U���u�u�u�9�2�}�W���Y���F�N��U����
�&�u�j�<�(���
����U��\�U���u�u�u�u�w�}������ƹF�N��U���=�;�4�
��.�Fہ�
����[�=N��U���u�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�0�|�#�8�}���Y���F�N��U���4�
��3�:�a�W���*����S��D��A�ߊu�u�u�u�w�}�W�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��A���8�d�n�u�w�}�W���Y����������u�u�u�u�w�5�Ͽ�&����GW��Q��D���k�_�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���PӒ��]l�N��U���u�u�u�u�w�<�(������F��h=����
�&�
�`�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�`�1�0�F��Y���F�N��U���;�u�3�_�w�}�W���Y�ƻ�V��G1��*���c�3�8�d�w�c�}���Y���F�N�����}�%�6�;�#�1����H����C9��G�����u�u�u�u�w�}�W���Y����C9��h��U��4�
��&�f�����O���F�N��U���u�0�&�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���O����lW��=N��U���u�u�u�u�w�3�W���s���F�N�����u�%��
�#�j����H���l�N��U���u�u�u�<�w�u��������\��h_��U���6�|�u�=�9�}�W���Y���F�N��U����
�&�u�j�<�(���
����U��Y�U���u�u�u�u�w�}����s���F�N��U���u�u�4�
��;���Y����g9��Y�����c�_�u�u�w�}�W���Y�Ʃ�WF��d��U���u�u�u�"�2�}����&����l ��h_�H���u�u�u�u�w�}�W������R��X ��*���<�
�u�u�'�>�^�����ƹF�N��U���u�u�u�u�'��(���Y����C9��h��L���8�d�n�u�w�}�W���Y�����Rd��U���u�u�u�u�w�}�WϿ�&����@�
N��*���&�d�
�&��j�}���Y���F�N�����<�n�u�u�w�}�W�������R��c1��Dӊ�&�
�m�h�w�}�W���Y���F���]´�
�:�&�
�8�4�(���Y����VO�C�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�e�1�0�F��Y���F�N��U���9�0�u�u�w�}�W���Y���F��G1��*���u�h�4�
��.�Fց�
����l�N��U���u�u�u�0�3�4�L���Y���F���ʴ�
��&�g��.�(��D��ƹF�N��U���u�u�3�}�6�����&����P9��
N��*���|�!�0�_�w�}�W���Y���F�N��*���3�8�i�u�'��(���H����lT��=N��U���u�u�u�u�w�1����Y���F�N��U���u�%��
�$�}�JϿ�&����GT��Q��D��u�u�u�u�w�}�W�������U]ǻN��U���u�u�=�;�6��#���K¹��^9��S����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�4�
��;���Y����g9��1����_�u�u�u�w�}�W���Y����9F�N��U���u�u�u�u�w�-�9���
�����d:�����3�8�g�n�w�}�W���Y���F��Y
���ߊu�u�u�u�w�}��������@F�NךU���u�u�u�u�w�}����&����[�o6��-���������/��Y���F��Y
�����_�u�u�;�w�/����B���F������u�&�<�;�'�2����Y��ƹF��G1�����&�<�;�%�8�}�W�������R��C��Yʴ�
�<�
�&�&��(���&����J��G1��Yʴ�
�<�
�&�&��(���H����lT��=N��U���<�_�u�u�w�}����Q������T�����2�6�d�h�6�����P�ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�����e�|�:�u��-��������Z��S�����|�4�1�}�'�>��������lW������6�0�
��$�o�(���&���O��_�����u�u�u�u�w�-����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�:�0�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�4�
�3�8�����Ƽ�\��D@��X���u�4�
�1�2�<����&����\��E�����%�&�4�!�w�-��������`2��C_�����|�u�u�7�0�3�W���Y����UF�Y��]���6�;�!�9�0�>�F������R��N�����%�6�;�!�;�:���DӇ��@��T��*���&�d�3�8�g�t�W������F�N��Uʴ�
�1�0�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��[��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������,�4�&�2�w�/����W���F�V�����
�&�<�;�'�2�W�������@N��h��U���&�2�6�0��	���&����V�N�����;�u�u�u�w�4�W�������]��[����h�4�
�0�w�3�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����ד�@��G��U���;�_�u�u�w�}�W���	����W�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�%�%�<���Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�u�u�6��������F��C1�����;�
�
�'�#���������T��h����u�%�'�!�%��W������C��R ��A���<�0�4�&�0����H¹��l�N��*��� �;�g�i�w�(�(�������lS��E��*���<�;�3�
�f�m���s���K��G1�����1�d�f�4�$�:�W�������K��N�����<�
�1�
�f���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����H���N��h�����#�
�u�u�'��(���Q�ƨ�D��_��N���u�0�1�%�8�8��Զs���K��G1�����1�d�`�4�$�:�W�������K��N�����<�
�1�
�d���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����J���N��h�����#�
�u�u�'��(���Q�ƨ�D��\��N���u�0�1�%�8�8��Զs���K��G1�����1�d�f�4�$�:�W�������K��N�����<�
�1�
�a���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����O���N��h�����#�
�u�u�'��(���Q�ƨ�D��X��N���u�0�1�%�8�8��Զs���K��G1�����1�d�f�4�$�:�W�������K��N�����<�
�1�
�`���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����N���N��h�����#�
�u�u�'��(���Q����\��XN�\��u�u�0�1�'�2����s���F������7�1�d�f�6�.��������@H�d��Uʴ�
�<�
�1��e�(�������A	��N�����&�4�
��1�0�}���Y����]l�N��U���u�u�u�4��4�(���&����[�V�����
�#�
�u�w�-�4���
������Y��D���n�u�u�0�3�-����
��ƓF�C�����2�7�1�g�a�<����Y����V��C�U���4�
�<�
�3��Fف�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F��*���&�
�#�
�w�}����&���� F��@ ��U���n�u�u�0�3�-����
��ƓF�C�����2�7�1�g�d�<����Y����V��C�U���4�
�<�
�3��E܁�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6��������� F�F��*���&�
�#�
�w�}����&����
F��@ ��U���n�u�u�0�3�-����
��ƓF�C�����2�7�1�g�g�<����Y����V��C�U���4�
�<�
�3��D߁�
����l��TN����0�&�4�
��;��ԜY�Ʈ�T��N��U���u�u�u�u�6���������F�F��*���&�
�#�
�w�}����&����U��X����|�n�u�u�2�9��������9l�N�U���&�2�7�1�e�j�����Ƽ�\��D@��X���u�4�
�<��9�(��&����T��E��Oʥ�:�0�&�4������s���Q��Yd��U���u�u�u�u�w�<�(���&����U��S�����:�&�
�#��}�W���:����^N��
�����d�|�n�u�w�8�Ϯ�����lǑN��X���%�&�2�7�3�o�BϿ�
����C��R��U���u�u�4�
�>�����Lƹ��@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9��N�U´�
�:�&�
�!��W���	����U��^�����:�g�|�n�w�}����	����@��=d��U���u�%�&�2�5�9�D���
������T��[���_�u�u�%�$�:����Jʹ��@��h����%�:�0�&�6��$������F��P��U���u�u�u�u�w�}��������W9��R��]����
�&�}�w�2����I���R��X ��*���
�|�_�u�w�3�W�������9lǻN��Xʴ�
�<�
�1��m�����Ƽ�\��D@��X���u�4�
�<��9�(�������]9��X��U���6�&�}�%������Y����V��=N��U���u�u�u�u�w�-��������F�F��*���&�
�#�
�w�}����&����F��@ ��U���n�u�u�0�3�-����
��ƓF�C�����2�7�1�c�w�.����	����@�CךU���%�&�2�7�3�k�(�������A	��N�����&�4�
��1�0�}���Y����]l�N��U���u�u�u�4��4�(���&���F��G1�����9�d�d�h�6��$�������W	��C��@���_�u�u�;�w�/����B��ƹF�N��*���
�1�
�l�6�.��������@H�d��Uʴ�
�<�
�1��d��������\������}�%��
�$�t�W�������9F�N��U���u�u�u�%�$�:����N���N��h�����#�
�u�u�'��(���Q�ƨ�D��V��N���u�0�1�%�8�8��Զs���K��G1�����1�m�d�4�$�:�W�������K��N�����<�
�1�
�b���������PF��G�����4�
��3�:�W�W�������F�N��U���u�u�4�
�>�����L���N��h�����#�
�u�u�'��(���Q�ƨ�D��Z��N���u�0�1�%�8�8��Զs���K��G1�����1�m�u�&�>�3�������KǻN�����2�7�1�m��.����	����	F��X��´�
��3�8�]�}�W������F�N��U���u�4�
�<��9�(��E����C9��Y�����d�h�4�
��;���Y����G	�G����u�;�u�'�4�.�L�ԶY���F��h��*���
�c�4�&�0�}����
���l�N��*���
�1�
�c�6�.���������T��]����
�&�|�w�}�������F�N��U���u�%�&�2�5�9�N���D�έ�l��D��ۊ�u�u�%���.�_������\F��G�U���0�1�%�:�2�.�}�ԜY�����D�����
��&�d��.�(���
������T��[���_�u�u�%�$�:����&����GW��Q��L���&�2�
�'�4�g��������C9��P1����f�_�u�u�2�4�}���Y���Z �V�����1�
�g�|�#�8�W���Y���F������6�0�
��$�l�(���&�����T�����2�6�d�_�w�}�W������F�N��U���4�
�<�
�$�,�$����֓�@��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����0�
��&�f�����HӇ��Z��G�����u�x�u�u�6�����
����g9��\�����d�4�&�2��/���	����@��G1�����1�m�|�u�w�?����Y���F��QN�����2�7�1�m�~�)����Y���F�N�����2�6�0�
��.�F݁�
����Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����9��Z1�U��4�
�:�&��2����B���F���U���u�u�u�0�3�-����
��ƓF�C�����2�6�0�
��.�F܁�
������^	�����0�&�u�x�w�}��������V��c1��Dي�&�
�g�4�$�:�(�������A	��D�����2�7�1�d�d�W�W�������F�N�����4�
�<�
�3��@�������9F�N��U���u�%�&�2�4�8�(���
����U��\��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-��������`2��C_�����d�u�h�4��2��������]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�%�&�2�4�8�(���
����U��]�����;�%�:�0�$�}�Z���YӇ��@��T��*���&�d�
�&��n��������\������}�%�&�2�5�9�E��s���Q��Yd��U���u�<�u�4��4�(���&������YNךU���u�u�u�u�'�.��������l��1����u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W���	����l��F1��*���a�3�8�d�w�`��������_	��T1����u�u�u�;�w�;�W���YӃ����T��N�ߠu�u�x�u�'�.��������l��1����u�&�<�;�'�2����Y��ƹF��G1�����0�
��&�f�����L����Z��G��U���'�6�&�}�'�.��������9F����ߊu�u�u�u�1�u��������lP�����ߊu�u�u�u�w�}��������B9��h��C���8�d�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƭ�l��h�����
�!�c�3�:�l�W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������B9��h��B���8�d�u�&�>�3�������KǻN�����2�6�0�
��.�F؁�
����l��^	�����u�u�'�6�$�u��������lT��d��Uʷ�2�;�u�u�w�}��������T9��S1�B���=�;�_�u�w�}�W���Y����Z��D��&���!�b�3�8�f�}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�j����H�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�l�3�8�f�}����Ӗ��P��N����u�%�&�2�4�8�(���
����U��V�����;�%�:�u�w�/����Q����Z��S
��C�ߊu�u�0�<�]�}�W���Y���R��^	�����c�u�=�;�]�}�W���Y���R��^	������
�!�l�1�0�F���DӇ��P	��C1�����d�_�u�u�w�}����s���F�N�����<�
�&�$����������F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��^	������
�!�
�$��W�������A	��D�X�ߊu�u�%�&�0�>����-����l ��h^�����;�%�:�u�w�/����Q����Z��S
��L�ߊu�u�0�<�]�}�W���Y���R��^	�����l�u�=�;�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�1��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�e�3�8�f�}����Ӗ��P��N����u�%�&�2�4�8�(���
����U��W�����;�%�:�u�w�/����Q����Z��S
��M���u�u�7�2�9�}�W���Yӏ����D�����d�f�u�=�9�W�W���Y���F��h��*���$��
�!�g�;���Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�<�
�&�&��(���I����lW��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h��*���$��
�!�f�;���Y����T��E�����x�_�u�u�'�.��������l��1����
�&�<�;�'�2�W�������@N��h��*���
�`�|�u�w�?����Y���F��QN�����2�7�1�g�b�}����s���F�N�����<�
�&�$����������F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�4�
�>�����*����W��D��E��u�%�6�;�#�1����I���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����<�
�&�$���݁�
����R��P �����&�{�x�_�w�}��������B9��h��*���
�
�&�<�9�-����Y����V��V�����1�
�d�|�w�}�������F���]���&�2�7�1�f�n�W������F�N��Uʴ�
�<�
�&�&��(���&����F������!�9�2�6�f�W�W���Y�Ʃ�@�N��U���u�u�4�
�>�����*����9��Z1�I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N��*���
�&�$���)�(���&�ƭ�@�������{�x�_�u�w�-��������`2��C]�����
�&�<�;�'�2�W�������@N��h��*���
�f�|�u�w�?����Y���F��QN�����2�7�1�d�b�}����s���F�N�����<�
�&�$���܁�
����[��G1�����9�2�6�d�]�}�W���Y����l�N��U���u�4�
�<��.����&����U��N�U���6�;�!�9�0�>�G�ԜY���F��SN��N�ߊu�u�;�u�%�>���s���K�V�����&�$��
�#�����Y����T��E�����x�_�u�u�'�.��������l��h��*ي�&�<�;�%�8�}�W�������R��^	�����d�|�u�u�5�:����Y����������7�1�g�c�w�5��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�d�_�w�}�W������F�N��U���4�
�<�
�$�,�$���ǹ��^9��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h��*���$��
�!��.�(���
������T��[���_�u�u�%�$�:����&����GS��D��*���<�;�%�:�w�}����
�έ�l��h��*���|�u�u�7�0�3�W���Y����UF��G1�����1�m�d�u�?�3�}���Y���F�V�����&�$��
�#�����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�<�
�&�&��(���&����F������!�9�2�6�g�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���R��^	������
�!�
�$��W�������A	��D�X�ߊu�u�%�&�0�>����-����l ��h[�����;�%�:�u�w�/����Q����Z��S
��E�ߊu�u�0�<�]�}�W���Y���R��^	�����e�u�=�;�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�1��ԜY���F�N��*���
�&�$���)�(���&�����T�����2�6�e�_�w�}�W����ƥ�FǻN�����'�6�&�n�]�}�W��Y����Z��D��&���!�
�&�
�w�.����	����@�CךU���%�&�2�6�2��#���N����lP��D�����:�u�u�'�4�.�_���
����W��]��U���7�2�;�u�w�}�WϷ�Yۇ��@��U
��D��u�=�;�_�w�}�W���Y�ƭ�l��h�����
�!�
�&��}�JϿ�&����G9��P��D�ߊu�u�u�u�;�8�}���Y���F�V�����&�$��
�#�����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����l��F1��*���
�&�
�u�$�4�Ϯ�����F�=N��U���&�2�6�0��	��������l��^	�����u�u�'�6�$�u��������lQ��=N��U���<�_�u�u�w�}����	����l��hY�U���;�_�u�u�w�}�W���	����l��F1��*���
�&�
�u�j�<�(���
����T��UךU���u�u�9�0�]�}�W���Y���R��^	������
�!�
�$��W������]��[����_�u�u�u�w�3�W���Y����������n�_�u�u�8�1����6����R��B1�@���u�h�}�8������K����]��E�� ��m�%�|�_�w�}��������F��X�� ��d�%�u�h��0�(������� V��V �����3�
�d�
�e�f�W�������K!��x��D���3�
�`�
�e�a�WǪ�	����U��W��Gʴ�1�2�%�3��l�(��B��� ��v,��:���d�f�3�
�d��F��Y����q5��B��@ي�0�
� �g�c�-�L���YӀ��r$��x��D���;�2�3�
�d��E��Yۏ��R
��V1�����;�
�0�
�e�o��������]��[�*��e�e�e�n�w�}����;����G9��1�����c�
�f�i�w�}�W���YӀ��r$��x��D���'�2�d�`�w�5��������l ��[�����|�h�r�r�w�1��ԜY���F��h/�����
�`�
�
�"�o�B���B��� ��v,��:���d�`�g�3��k�(��E�ƪ�l'��O!��*���
�0�
� �e�m���Y����`9��d����`�g�!�
�9����I����[��d1��&���!�d�`�'�0�l�B��Y����`9��d����`�3�
�e��m�K�������R9��=N��U������!�f�h����I����Z�V�����
�#�g�f�f��G��Y����`9��d����`�;�2�3��k�(��E����`9��d����`�g�!�
�9�����K����\��G1�����9�f�
�e�g�m�G��Y����`9��d�����!�
�;�
�"�o�B���Y����`9��d����`�d�3�
�a��D�ԜY�ƪ�l'��O!��*��� �g�f�%�w�`�}���Y���Z��[��*���=�;�}�8�����I����O�I�\ʰ�&�u�u�u�w�}����;����G9��1��*��
�d�_�u�w��6���6����\9��C1��*��
�d�i�u���$�������F9��1��N���u�3�
�!�f�o�E���&����CU�
NךU���u�u�;�4�'�<�Fϩ�����V
��Z�����g�
�g�e�w�}�F�������9F�N��U���6�
�d�
�"�h�@���B��� ��T��D؊�
� �`�d�'�}�J�ԜY���F��h/�����
�`�
�
�"�o�B���Y����N��[1��݊� �a�`�%��t�J���^�Ʃ�@�N��U���3�
�!�d�e�o����Lǹ��l�N��*���d�g�a�3��j�(��E��ƹF�N��&�����!�d�b�/���L�ƻ�V�D�����
� �`�`�'�u�^��^���V
��d��U���u�3�
�!�f�o�B���&����CU��N�����!�d�g�`�1��Aց�J���9F�N��U������!�f�n����Jʹ����YN�����8�f�3�
�o��E��Y���O��[�����u�u�u��4��F݁�&����W��UךU����6�
�d��(�B���	���l�N��Uʼ�
�9�=�
�w�5��������F9��1��]���h�r�r�u�;�8�}���Y���U5��u=�� ���`�
� �g�n�-�L���YӀ��P��W��*���`�`�%�u�j�W�W���Y�ƪ�l'��O!��*���
�0�
�g�`�*����
����^��Q��@ߊ�g�e�u�u�f�t����Y���F������d�
� �`�o�-�L���YӀ��P��W��*���`�g�%�u�j�W�W���Y�ƪ�l'��O!��*���
�0�
�g�`�*����
����^��Q��Mڊ�g�e�u�u�f�t����Y���F������d�
�
� �b�h���Y����`9��h_�*ފ� �c�a�%�w�`�}���Y���U5��u=�� ���`�
�0�
�e�j� ���Yە��l��1��*��
�g�e�u�w�l�^ϻ�
��ƹF�N��&���
�d�
�
�"�k�A���B��� ��T��Dӊ�
� �`�l�'�}�J�ԜY���F��h/�����
�`�
�
�"�o�B���Y����N��[1��Ҋ� �`�`�%��t�J���^�Ʃ�@�N��U���3�
�!�d�n�n����J����l�N��*���d�l�c�3��e�(��E��ƹF�N��&�����!�d�b�o����Oƹ����YN�����3�
�b�
�e�m�W���H����_��=N��U���u�����)�F�������S��=N��U���6�
�d�
��(�B���	���l�N��Uʳ�
��-� ��h�(���&������YN�����8�g�3�
�e��E��Y���O��[�����u�u�u��4��Fց�&����R��UךU����6�
�d�����A����[�N��U���3�
��-�"��Bځ�&����S��N�����&�9�!�%��(�C���	����[�I�����u�u�u�u�w�;�(���H�ߓ�l ��W����u�u�3�
�#�l�N�������9��R�����u�u�u����8���H�ӓ�l ��X�����=�;�}�0��0�D���&����CT�N��R��u�9�0�_�w�}�W���*����W��1��*��
�f�_�u�w�����Hʹ��lS��h�I���u�u�u�u�1��5�������9��P1�@���=�;�}�0��0�E���&����CT�N��R��u�9�0�_�w�}�W���*����K)��h_�*؊� �g�`�%�l�}�Wϸ�&����9��Q��Eӊ�f�i�u�u�w�}�Wϸ�&����|��[�����f�
�d�"�2�}����&����_��F�U���d�|�0�&�w�}�W���YӀ��r$��x��D���g�3�
�c��l�}���Y����G9��h\�� ��l�%�u�h�]�}�W���Y����q5��B��@ي� �g�l�%�w�5��������CT��B1�F���}�|�h�r�p�}����s���F�Q=����
�
� �a�n�-�L���YӀ��P��1�����c�
�f�i�w�}�W���Yӏ��R
��V1����u�&�9�!�'����L����O�I�\ʰ�&�u�u�u�w�}��������9��hZ�*��_�u�u��4��O�������9��R�����u�u�u�;�6�-���������h��M���
�e�
�g�g�}�W��PӃ��VFǻN��U����6�
�m�b�;�(��&����F�Q=����
�
� �a�a�-�W��s���F�Q=��7��� �
�`�
�2��E��������h��F���
�m�
�g�g�}�W��PӃ��VFǻN��U����6�
�m�d�;�(��&����F�Q=�����&�
�!� �#�/�(���K����_��G]��H�ߊu�u�u�u�2��C������G��D1����d�}�|�h�p�z�W������F�N��*����g��!�f�l�D�������
]ǻN��&���
�4�0��%�>����M¹��U��Y��F��u�u�u�u�w�;�(���5�Ԣ�F��_��*���
�f�l�"�2�}��������l��h_�M��u�u�d�|�2�.�W���Y��� ��T������'�6� �2�i�(���@�֓� ]ǻN��&���
�4�0��%�>����M¹��U��]��F��u�u�u�u�w�/���Jӑ��]F��R����
�0�
�f�b�m�W���H����_��=N��U���u��6�
�6�8�$�������lR��1��*��
�f�_�u�w���������G��C��*���l�3�
�f��n�K���Y���F��R	��A���=�;�}�0��0�Fց�����T�N��R��u�9�0�_�w�}�W���*����p��h=�� ���'�
�d�`�1��E܁�J���F��h��6���
�!� �!�%��F���&����CU�
NךU���u�u�0�
�c�}����Q����\��h��*��d�e�u�u�f�t����Y���F������4�0��'�4�(���&����l^��h����u��6�
�6�8�$�������lR��1��*��
�f�i�u�w�}�W�������f*��Y!��*��
�
�0�
�d�d� ���Yۉ��P	��1����a�}�|�h�p�z�W������F�N��*����&�
�!�"�)����A����_��G]�U���3�
�!��$���������^��h��L���%�u�h�_�w�}�W������� F��R �����!�%�`�'�0�l�C���P���A�R��U���u�u�u�3��)�4���&����P��R1�*ۊ� �l�m�%�l�}�Wϸ�&����R��d�����0�a�
�
�"�d�F���Y���F�N�����d�l�"�0�w�.����	�ѓ�V��[�E���u�d�|�0�$�}�W���Y����`9��h-�����'�6� �0�c��(���@�ғ� ]ǻN��&���
�4�0��%�>����M˹��U��V��F��u�u�u�u�w�;�(���5�Ԣ�F��_��*���
�f�l�"�2�}��������l��h_�G��u�u�d�|�2�.�W���Y��� ��T������'�6� �2�i�(܁�����l��=N��U���6�
�4�0��/��������U��Y��F��u�u�u�u�w�/���Jӑ��]F��Z��*���
�f�a�e�w�}�F�������9F�N��U���
�a�n�u�w�;�(���:����`��T�����
�
� �l�b�-�W��s���F�E��D��"�0�u�:��2�ށ�����W�N��R��u�9�0�_�w�}�W���*����p��h=�� ���'�
�`�3��m�(��s���U5��C1�����!� �!�'��h�E���&����CU�
NךU���u�u�0�
�c�}����Q����G��1����a�}�|�h�p�z�W������F�N��*����&�
�!�"�)����L�ד�F9��1��N���u�3�
�!��.�(�������V9��h]�� ��l�%�u�h�]�}�W���Y����~3�� ����d�f�'�2�f�j�W����ο�_9��G_�����d�`�}�|�j�z�P������F�N�����!��&�
�#�(����&�ӓ�l ��Y����u�u�3�
�#���������F��[��*���l�`�%�u�j�W�W���Y�ƾ�T9��N�����&�9�!�%�n�/���O����[�I�����u�u�u�u�w�;�(���:����`��T�����
�
� �l�n�-�L���YӀ��P��V��&���6� �0�`��(�N���	���l�N��Uʳ�
���g��)�F���J����lW��N�����!�%�&�'�0�l�F���P���A�R��U���u�u�u�'�0�l�D�ԜY�ƪ�l��Z_�����;�0�4�1��8����&¹��lW��1��U��_�u�u�u�w�-��������9��@��U²�%�3�
�f��o�G���Y�����RNךU���u�u��6��<��������A��1�����d�e�n�u�w�;�(���¹��l4��P�����:�'�0�c�1��F���	���l�N��Uʴ�
�:�&�
�!�o�Gϩ�����A��B1�F���}�|�h�r�p�}����s���F�Q=�����&�
�!� �#�/�(���@����lW��UךU����!�'�d������&����p	��T��*���d�b�
�f�k�}�W���Y����C9��Y����
�u�=�;��/�(���H�ޓ�N��S��D���0�&�u�u�w�}�Wϸ�&����R��d�����0�a�
�
�2��D��s���U5��v*��:����1�d�c�1��Gށ�H���A��Z����u��-� ��3����O¹��U��]��F��u�u�u�u�w�;�(���5�Ԣ�F��_�� ��d�%�u�=�9�u��������U�� Y��G��u�u�d�|�2�.�W���Y�����h_�N���u�3�
���o�8���H�ד�F9��1��U��%��&�9��l����Mʹ��l�N��*����g��!�f�l��������9��hY�*��i�u�!�
�8�4�(�������]��Y�����&�9�
�
�"�j�F���P����]��Y�����:�&�
�#�c�n�1���?���l�N��*����g��!�f�l����	����l �� Y�����h�_�u�u�w�}����&����P��h�����
�a�
�f� �8�Wǭ�����V��B1�B���}�|�h�r�p�}����s���F�D�����
� �b�f�'�f�}���Y����A��B1�M���6�1�u�&�>�3�������KǻN����� �d�m�:�4�9�(�������A	��N�����&�4�
�<��.����&����U��B�����2�6�0�
��.�D������R��^	������
�!�e�1�0�F��
����^��1�����4�
�0�
�c�e�W���
����@��d:�����3�8�g�|�w�}�������F���]���%�6�;�!�;�:���DӇ��@��T��*���&�g�
�&��m�W���Yە��l��X�����'�4�
�0��i�O������]��[��E���u�=�;�_�w�}�W���Y�ƫ�C9��h_�*���:�0�i�u�'�>�����ӓ�l�N��Uʰ�&�3�}�}�'�>��������lW������6�0�
��$�n����K�ƣ�N��h�����:�<�
�u�w�-��������`2��C\�����d�|�|�!�2�}�W���Y���F��E�� ��m�:�6�1�w�`��������_��UךU���u�u�9�<�w�u��������\��h_��U���&�2�6�0��	��������O��_�����u�u�u�u�w�/�(���H�ޓ�C��RN�U���6�;�!�9�b�o�}���Y���V
��d��U���u�u�u�2�'�;�(��&����W�
N��-���w�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����^��N�����u�'�6�&�y�p�}���Y����U��V��E���&�2�
�'�4�g��������]9��G��D���%�&�2�6�2��#���K����lW�V�����&�$��
�#�����UӀ��P��V��&���6� �0�a�����I���� ��T������'�6� �2�i�(ց�����
V�V�����&�$��
�#�m����H����C9��P1������&�g�
�$��G�ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��G1�����0�
��&�e�����I����[��=N��U���u�u�u�'��(�F���	��� ��T������'�6� �2�i�(ց�����
V��N��U���0�&�3�}�6�����&����P9��
N��*���
�&�$���)�G�������F��R ��U���u�u�u�u�0�-����I˹��Z�Q=�����&�
�!� �#�/�(���@����
U��G]�U���u�u�0�&�1�u�_�������l
��^��U���%�&�2�6�2��#���K����lW�X�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�~�)����Y���F�N����� �d�m�%�w�`��������]ǻN��U���9�0�_�u�w�}�W���Y����U��V��E��u������/���!����k>��o6��-����n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϹ�	����V��G_�����;�%�:�0�$�}�Z���YӁ��l ��^��ۊ�&�<�;�%�8�}�W�������R��^	������
�!�
�$��[Ͽ�&����P��h=�����3�8�g�u�'�.��������l��1����y�4�
�<��.����&����l ��h\����u�0�<�_�w�}�W�������C9��Y�����6�d�h�4��4�(�������@��h��*��|�!�0�u�w�}�W���Y����A��B1�M���u�h�4�
�8�.�(���K�Պ�V��UךU���u�u�9�<�w�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��EN�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�g�u�%�u��������\��h_��U���&�2�6�0��	���&����V�N�����u�u�u�u�w�}��������9��R�����:�&�
�#�e�m�}���Y���V
��d��U���u�u�u�2�'�;�(��&���F��o6��-���������/���!����k>�=N��U���u�;�u�3�w�}�Wϻ�Ӗ��P��dװU���x�u�'�
�"�l�C�������R��P �����&�{�x�_�w�}��������l	��X
�����2�
�'�6�m�-����
ۇ��@��T��*���&�g�3�8�f�}��������B9��h��*���
�y�4�
�>�����*����V��D��L���0�
�8�d�a�9��������T9��]����<�
�&�$����������OǻN�����_�u�u�u�w�;�_���	����@��X	��*���u�%�&�2�4�8�(���
����U��^�����}�0�
�8�f�k��������A��Z�U���%�6�;�!�;�l�G���Y����l�N��U���u�2�%�3��l�(������F��h�����#�
�n�u�w�}�Wϻ�
���N��h�����:�<�
�u�w�-��������`2��C]�����|�:�u�4��2��������F�V�����&�$��
�#�m����H�����YNךU���u�u�u�u�%����M����\��S�����;�!�9�`�d�W�W���Y�Ʃ�@��F��*���&�
�:�<��}�W���
����@��d:��؊�&�
�|�u�?�3�}���Y���F�P�����d�
�%�:�2�a�W�������l
��h\�U���u�u�0�&�w�}�W���Y�����h��D���:�6�1�u�j��/���[���F�N��ʼ�n�_�u�u�9�}����
��Ɠ9F�C����3�
�d�
�g�<����Y����V��C�U���2�%�3�
�f��G���
����C��T�����&�}�������L����lW�� B�����2�6�0�
��.�E������R��^	������
�!�
�$��[Ͽ�&����P��h=����
�&�
�l�w���������G��C��*���l�3�
�`��n�W�������@��C�����
�m�l�'�0�l�N������T9��R��!���g�
�&�
�g�W�W�������F�N�����}�%�6�;�#�1����H����C9��P1������&�g�
�$��G�������9F�N��U���u�'�
� �f�i����DӀ��P��V��&���6� �0�a������J����F�N�����3�}�4�
�8�.�(�������F��h��*���$��
�!�g�;���P�Ƹ�V�N��U���u�u�2�%�1��Fہ�I���U5��C1�����!� �!�'��e�N���&����CU��N��U���0�&�3�}��-��������Z��S�����2�6�0�
��.�E������\�V�����
�:�<�
�w�}��������B9��h��*���
�|�|�!�2�}�W���Y���F��E�� ��a�%�u�h�1��5�������9��P1�@��u�u�u�u�2�.�W���Y���F�	��*���d�a�%�u�j��/���!����k>��o6��-���������}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��G1��*��
�d�4�&�0�}����
���l�N�����
�d�
�d�6�.���������T��]���&�2�6�0��	��������F��h��*���$��
�!��.�(������T9��R��!���g�
�&�
�n�}��������B9��h��D���8�g�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���e�3�8�d�~�}����s���F�N�����3�
�d�
�f�a�W�������l
��1��M��e�n�u�u�w�}�������R��X ��*���<�
�u�u�'�.��������l��h��*���:�u�4�
�8�.�(�������F��h��*���$��
�!��.�(�������C9��Y�����6�d�h�4��4�(�������@��h��*��|�u�=�;�]�}�W���Y���T��Q��Dފ�d�i�u�%�4�3����J����9F�N��U���0�_�u�u�w�}�W�������lW��h�I���������/���!����k>��o6��-���n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������
9��T��U���<�;�%�:�2�.�W��Y����A��B1�L���6�1�
�&�>�3����Y�Ƽ�\��DF��*���
�&�$���)�(���&����C9��P1������&�g�
�$��N�������CW��h
�����;�'�2�d�c�q��������V��c1��Gۊ�&�
�e�_�w�}����s���F�^��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�d�3�8�e�t����Q����G��X�����2�;�'�2�f�i�W���	����@��A_��\���!�0�u�u�w�}�W���YӁ��l ��_�����1�u�h�4��2����ƹ��9F�N��U���<�u�}�4��2��������F�V�����&�$��
�#�����PӉ����T�����2�6�d�h�6�����
����g9��^�����l�|�u�=�9�W�W���Y���F��G1��*��
�%�:�0�k�}��������ES��d��U���u�0�&�u�w�}�W���Y����A��B1�L���6�1�u�h�u��/���s���F�R ����_�u�u�;�w�/����B��ƹF�N�����
�d�
�e�6�.��������@H�d��Uʲ�%�3�
�d��m��������\������}�%�&�2�4�8�(���
�Փ�@��N��*���
�&�$���)�G������� ��T������'�6� �2�h�(ׁ�����l�������4�0��'�4�(���&˹��T9��\����<�
�&�$����������J��d1��&���!�&�3�
�c��D�ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��G1�����0�
��&�e�����I����[��=N��U���u�u�u�'��(�F���	��� ��T������'�6� �2�h�(ׁ�����T��N��U���0�&�3�}�6�����&����P9��
N��*���
�&�$���)�G�������F��R ��U���u�u�u�u�0�-����Hʹ��Z�Q=�����&�
�!� �#�/�(���A����
^��G]�U���u�u�0�&�1�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O�C��U���u�u�u�u�w�:����&����CV�
N��*���-� �
�
�"�o�D���B���F����ߊu�u�u�u�w�}��������l��S��-���������/���!����k>��o6��N���u�u�u�0�3�4�L�ԜY�Ʃ�WF��X���ߠ_�u�u�x�0�-����Hʹ����^	�����0�&�u�x�w�}��������
9��h�����%�:�u�u�%�>����	����l��F1��*���
�&�
�y�6�����
����g9��^�����l�u�%�&�0�>����-����9��Z1�Yʳ�
��-� ��h�(ށ�����l��=N��U���<�_�u�u�w�}��������]��[����h�4�
�<��.����&����l ��h\�\ʡ�0�u�u�u�w�}�W�������F9��1��U��4�
�:�&��+�E��s���F�R�����4�
�:�&��2����Y�ƭ�l��h�����
�!�e�3�:�l�^������F�N��U���2�%�3�
�f��F��Y����\��h��G���m�e�e�n�w�}�W�������N��G1�����9�2�6�d�j�<�(���&����l5��D�����g�|�!�0�w�}�W���Y�����h��D���%�u�h�3������&����9��h\�*��_�u�u�u�w�1��ԜY���F�N�����
�d�
�d�k�}�/���!����k>��o6��-���������L���Y�������U���u�0�1�%�8�8��Զs���K��E�� ��m�%�u�&�>�3�������KǻN����� �d�m�%��.����	����	F��X��´�
�<�
�&�&��(���I����lW����*���3�
�e�d�'�q����J����T9��]����<�
�&�$����������OǻN�����_�u�u�u�w�;�_ǿ�&����G9��P��D��4�
�<�
�$�,�$����ד�@��G�����u�u�u�u�w�}�WϹ�	����T��G^��Hʡ�%�f�
�0��i�D�ԜY���F��D��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�e�3�8�f�t�W������F�N��Uʲ�%�3�
�g��m�K�������l ��^�*��_�u�u�u�w�1��ԜY���F�N�����
�g�
�e�k�}�/��Y���F��Y
�����u�u�0�1�'�2����s�����h��D���%�u�h�}�%����A����R��P�����e�
�g�n�]�}�W������F9��1��U���<�;�%�:�2�.�W��Y����A��B1�F���
�&�<�;�'�2�W�������@N��h��*���$��
�!�g�;���UӒ��lU��Q��D���%�y�!�%�d�����M���R��^	������
�!�d�1�0�E���Y����V��=N��U���u�3�}�4��2��������F�V�����&�$��
�#�l����K���G��d��U���u�u�u�2�'�;�(��&���F��G1�*���
�a�m�_�w�}�W�������N��h�����:�<�
�u�w�-��������`2��C\�����d�|�u�=�9�W�W���Y���F��G1��*��
�e�i�u�:��O���&����l��=N��U���u�9�0�_�w�}�W���Y�ƫ�C9��h_�*��i�u��n�w�}�W�������U]�N�����%�:�0�&�]�}�WϹ�	����U��G\��H���'�
� �d�d�-�W���Y����U��Z��G��_�u�u�x�0�-����J˹����^	�����0�&�u�x�w�}��������9��h�����%�:�u�u�%�>����	����l��F1��*���e�3�8�d�{�)���&����P��G\����a�
�0�
�c�n�W���
����@��d:�����3�8�g�|�w�}�������F���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�d�3�8�e�t�W������F�N��Uʲ�%�3�
�f��m�K�������l��h_�F�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
����U��W��U���;�_�u�u�w�}�W�������lW��h�I���8�
�f�3��l�D���B���F����ߊu�u�u�u�w�}��������l��S��-��u�u�u�u�2�9���s���V��G�����_�u�u�2�'�;�(��&���F��E�� ��m�%�u�;�w�/�(���H�ߓ�O��=N��U���2�%�3�
�d�>�W�������A	��D�X�ߊu�u�'�
�"�d�(�������]9��X��U���6�&�}�%�$�:����&����GW��D��Yʴ�
�0�u�%�$�:����&����GT��D��Yʴ�
�<�
�&�&��(���&����J��G1�����0�
��&�f�����K�ƭ�l��h�����
�!�e�3�:�l�[Ͽ�&����P��h=����
�&�
�e�]�}�W������F�N��U���4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t��������C9��Y�����6�d�h�4��8�^ϱ�Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���}�%�6�;�#�1����H����C9��P1������&�f�3�:�o�W���Q����\��h�����u�u�%�&�0�>����-���� 9��Z1�\ʺ�u�4�
�:�$�����&���R��^	������
�!�e�1�0�F�������C9��Y�����6�d�h�4��4�(�������@��h��*��|�u�=�;�]�}�W���Y���T��Q��F���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W�������l_��T��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F�	��*���l�
�e�4�$�:�W�������K��N�����3�
�f�%��.����	����	F��X��§�2�d�f�u�2��C������l_��1����g�y�4�
�>�����*����9��Z1�U���-� ��;�"��Aށ�&����U��N��*���
�&�$���)�(���&����C9��P1������&�d�
�$��[Ͽ�&����P��h=����
�&�
�f�w�-��������`2��C_�����d�|�u�u�5�:����Y�����F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�5��ԜY���F�N�����
�f�%�u�j�;�(���5�Ԣ�F��_��*���
�f�l�_�w�}�W�������N��h�����:�<�
�u�w�-��������`2��C_�����l�|�!�0�w�}�W���Y�����h��Lي�e�i�u�0��i�L���Y�����^��]´�
�:�&�
�8�4�(���Y����Z��D��&���!�
�&�
�~�2�Wǿ�&����G9��P��D��4�
�<�
�$�,�$����ѓ�@��G��U���;�_�u�u�w�}�W�������l_��G^��Hʧ�2�d�f�_�w�}�W�������N��h�����:�<�
�u�w�-��������`2��CZ�����|�u�=�;�]�}�W���Y���T��Q��F���u�h�3�
�#�d�(ہ�����W��N��U���0�&�u�u�w�}�W���YӁ��l ��]��E��u������/���!����k>��o6��-����n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϹ�	����
U��N�����u�'�6�&�y�p�}���Y����U��1��*���<�;�%�:�w�}����
�Υ�l��h\����d�f�u��4��Fց�&����U��N��*�����!�d�`�/���O����C9��P1������&�b�3�:�k�W���
����@��d:��ފ�&�
�y�4��4�(�������@��h��*���4�
�<�
�$�,�$����ғ�@��B�����2�6�0�
��.�F؁�
����l�N�����u�u�u�u�>�}�_�������l
��^��U���%�&�2�6�2��#���Hǹ��^9��G�����_�u�u�u�w�}�W���&���� 9��R�����d�f�_�u�w�}�W��������T�����2�6�d�h�6�����
����g9��^�����|�:�u�4��2��������F�V�����&�$��
�#�j����H�����YNךU���u�u�u�u�%����&���F��h��1���!�d�b�'�0�l�A��Y���F��[��U���%�6�;�!�;�:���DӇ��@��T��*���&�b�3�8�a�t����Y���F�N��U���
� �l�
�f�a�W�������l�N��Uʰ�&�3�}�4��2��������F�V�����&�$��
�#�����P�Ƹ�V�N��U���u�u�2�%�1��D���Y����`9��h_�*ߊ�0�
�f�c�]�}�W���Y����l�N��U���u�2�%�3��n����D�Ĕ�k>��o6��-���������/���!����F�N�����<�n�_�u�w�3�W�������9lǻN��Xʲ�%�3�
�b�4�}����Ӗ��P��N����u�'�
� �n�����
����C��T�����&�}�%�6�{�<�(���&����l5��D�����`�u�%�&�0�>����-����l ��h]����<�
�&�$���ځ�
����9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������_	��T1�Hʴ�
�<�
�&�&��(���&����O��EN�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�f�u�%�u��������\��h_��U���&�2�6�0��	��������O����ߊu�u�u�u�w�}��������P�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�'��(�N؁����R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�w�}��������l��S��&���
�d�
�
�2��D��s���T��Q��B���u�h�3�
�#�l�N������� U��=N��U���%�
� �c�n�-�W��[����[����*���3�
�g�
�d�`��������_��G�����w�w�_�u�w�>�؁�����lP��h�I���<�8�b�3��o�(������C9��Y�����d�n�u�u�>�0�(���J�ߓ�F�L�U���;�}�8�
�`�;�(��&�����T�����g�e�u�9�2��U�ԜY�ƥ�^��X�� ��f�%�u�h��>����&����CT��X�����;�!�9�d�f�f�W�������C��1��*���
� �d�a�'�}�JϷ�&����R9��=N��U���
�
�
� �`�h����DӀ��K'��N!��*���
�b�
� �`�l����J�����Y��E��u�u�9�6��o����@Ĺ��Z�G1��؊�
� �l�f�'�u�GϺ�����U�=N��U���
�
�
� �f�m�(��E�Ƽ�e��h_�� ��f�%�}�f�z�l��������l�N�����a�3�
�e�o�-�W��	����9��Q��E���%�}�e�1� �)�W��B���
��h8��*���d�c�
�d�k�}�(���K�ԓ�F9��Z��D��u�u�u�:�9�2�G��Y����\��hX�� ��d�
�a�i�w�����J����W��h�F���:�;�:�g�~�W�W�������9��h_�L���u�h�%��;��(���H����CW�N�Dʱ�"�!�u�|�]�}�W���&����lQ��h�I����-��,�"�����NŹ��lQ��h�F���:�;�:�g�~�W�W�������9��h_�D���u�h�w�w� �8�Wǲ�����l ��_�*��h�4�
�:�$��ׁ�?�Ʃ�@�L�U���;�!�=�g�1��G؁�K���V�@��U¡�%�d�
� �f�n����Y����\��h��*���u�9�0�w�u�W�W�������9��h]�*��i�u�e�u�?�3�_���&�ߓ�F9��1��U���%�6�;�!�;�e�1�������W�=N��U���9�&�
� �d�l����D������YN�����d�3�
�l��i�JϿ�&����G9��1��\ʰ�&�u�d�n�w�}�����Г�F9��W��G��u�e�u�=�9�u����&����l_��h�Hʴ�
�:�&�
�!��1������D��N�����=�m�3�
�g�m����D������YN�����
�
� �d�b��C������]��[��3���0�&�u�d�l�}�Wϰ�����U�� \��G��u�e�u�=�9�u��������l��
N��*���&�
�#�
��}����[����F�Y�����3�
�d�b�'�}�J���[ӑ��]F��X��*݊� �d�g�
�f�`��������_��h^�����u�e�n�u�w�3����K����W��G\��H���w�"�0�u�#�-�F܁�����l��
N��*���&�
�#�f�g�}����[����F�Y�����3�
�d�
�e�a�W��Y����N��G1�*���g�d�%�u�w�-�������� 9�������w�_�u�u�8�/�ځ�����l��S��D���=�;�}�8��o����Iʹ��[��G1�����9�g�
�|�2�.�W��B�����E��*���d�f�
�g�k�}�F������_	��a1�����e�b�%�u�w�-�������� 9�������w�_�u�u�8�/�ׁ�����9��R��W���"�0�u�9�4��B���&����l��
N��*���&�
�#�f�g�}����[����F�Y����� �d�m�%�w�`�U���������h_�� ��m�%�u�u�'�>��������O��[��W���_�u�u�'�4�3�F���&����CT�
N�����
� �c�l�'�}��������lU��h�N���u�:�!� �2�>����&����V9��D��*���d�f�
�f�k�}�W���Y����V
��Z�*���d�g�
�f� �8�Wǭ�����^��S�����
�0�
�a�o�m�W���H����_��=N��U���u��!�'�f��(�������W9��R��*܊�
� �d�d��n�}���Y����e��T��*ފ�'�!�
�&�>�3����K�ד� F�d��U���u�&�9�!�'�l����K�ғ� F��R �����!�%�b�
�2�2��������U��G��U��|�0�&�u�w�}�W�������A��~ �����
�;�
�:�%�8�A���&����l��=N��U���
�%�'�0�#�h� �������Z��Q��D���%�u�h�_�w�}�W�������CT��Q��D���%�u�=�;��8�(���H�Г�V��P�����d�d�}�|�j�z�P������F�N�����0�8�
�;��3��������A�� 1��*��c�%�n�u�w�-�G��&¹��l^��h�I���u�u�u�u�6�����&����lV��_��]���
�m�3�
�g��E��Y���O��[�����u�u�u�:���(���N�ӓ�]ǻN��*��� �!�d�
�"�e�N���Y���U5��v*��:����1�d�c�1��Gށ�H����W	��C��D���u�8�
�b�1��Cށ�J��ƹF��h<�� ���&�3�
�m��n�K�������]��[�*���u�:�
�
�"�j�B���P���F��a��*ۊ� �l�f�%�w�`��������V9��E�� ���a�
�
� �n�m���Y����l0��1�����e�a�%�u�j�;�(���:����`��T����
�
� �l�o�-�L���YӖ��R
��1��*��`�%�u�h�1�����
����A��B��@ߊ�
� �l�`�'�f�W�������l��h�����&�
� �b�b�-�W��s���F�V�����
�#�`�`�g�*��������l��1��*��
�g�e�u�w�l�^ϻ�
��ƹF�N�����;�!�9�d��m�L���YӔ��l��h��B���%�u�h�_�w�}�W���	����@��A_��A��u�=�;�}�:��(���J����T��G\��\��r�r�u�9�2�W�W���Y�ƭ�l��D�����a�e�n�u�w�/����&����CT�
N�����-���!�f�m����Lƹ���������!�9�d�d�l�}�Wϭ�����V��B1�B���u�h�}�8��d��������
9����U���
�8�l�3��k�(��B�����h��D���1�8�'�4��(�A���	���N��h��ۊ� �c�`�%�w�/����H����lP��h�N���u�&�9�!�'�l����Oƹ��Z�_�����u�3�
���o�8���H�ד�]9��c��*���b�f�%�u�w�-��������9��^�����u�e�n�u�w�.����	����W��E	��*���c�f�%�u�j�u��������l��X�����
�c�
�g�8�}����&����
W��G�U���&�9�!�%�e�;�(��&���F�N�����3�
���e����H����U��G�� ��f�%�u�u�'�>��������V�������w�_�u�u�2����&����A��h��A���%�u�h�}�2���������T��Q��F݊�g�:�u�8�����H����l�N�����%�f�3�
�`��E��Yە��l��_�� ��`�%�u�'�$�1����K����Q��G\����u�0�
�8�f����J����[�U��*���,� �
�`��(�D���	�ƣ���GY����� �c�b�%�~�W�W�������CW��Q��@ӊ�g�i�u�!�'�l�(���O�ד�F��SN�����%�a�3�
�b��E��Y����V
��Z�C���8�'�4�
�"�l�Cׁ�K�����h��D���%�u�'�!�'�l�(�������l ��^�*��n�u�u�&�;�)��������9��R��]���
�8�d�c�3�0����&����S��N��ʴ�
�:�&�
�!��^�ԜY�ƿ�_9��G_�*���:�2�;�3��l�N���Y���T��Q��Fي�g�:�u�8��h��������U��V�����_�u�u�0��0�F؁�����l��S�����m�3�
�l��o����
����^��h��C���%�|�_�u�w�8�(���H�Г�V��P�����d�e�%�u�j�u��������l��X�����f�1�8�'�6����Mƹ��]ǻN�����8�d�
� �a�d����D�ο�_9��G_�*���:�2�;�3��e�(������C9��Y�����d�n�u�u�$�1����@����_��G\��H���8�
�
� �d�j�����ƿ�_9��G_�����m�
�g�n�w�}��������U��Y��G��u�<�8�
�"�n�N���Y����R��X ��*���
�|�_�u�w�8�(���Kù��lW��1��U��_�u�u�u�w�-��������9��t^�E���=�;�}�8��j��������A��Z�]���h�r�r�u�;�8�}���Y���R��X ��*���g�f�m�e�g�f�W���
����^��h��D��
�f�i�u�w�}�W�������]��[�*ݓ�e�e�e�"�2�}����Kƹ��^	��V �����a�f�e�u�w�l�^ϻ�
��ƹF�N�����;�!�9�f���G��I���F��[1�����1�8�'�4��(�C���	���N��[1�����1�8�'�4��(�C���	�ƣ���hW�� ��b�%�|�_�w�}��������U��\�����h�_�u�u�w�}��������EU�� (��E��u�=�;�}�:��D�������]9��P1�F���|�h�r�r�w�1��ԜY���F��h�����#�g�f�m�g�m�L���Yӕ��l��1��*��
�g�i�u�%�+����Aƹ������*���d�3�
�d��o�L���Yӕ��l��1��*��
�g�i�u�#�-�N���&����CT��Y
�����8�
� �a�c�-�^�ԜY�ƿ�_9��GZ�� ��f�%�u�h�]�}�W���Y����Z9��Q��Fۊ�f�"�0�u�#�-��������
9��^��H��r�u�9�0�]�}�W���Y����\��h��@��e�_�u�u�2���������
9��R��]���
�8�g�
�2�2�������� 9����U���6�;�!�9�f�l�L���Yӕ��l��1�����4�
� �a�`�-�W��Q����l ��Y�����'�'�#�3��e�(��B�����h��C���
�a�
�g�k�}����&����|��[�����`�
�g�4�3�4��������lR��h�N���u�&�9�!�'����L����[�C��M���
�l�
�g�6�9��������U��W��G��u�u�&�9�#�-�(���L�ӓ�F�F�����3�
�e�
�e�<�ϭ�����9��hZ�*��n�u�u�&�;�)�ց�����l��S�����<�<�3�
�f��EϦ�Ӈ��P	��C1��D��n�u�u�&�;�)����&����CT�
N�����8�d�
�0�8�:����&����CT��X�����;�!�9�d�f�f�W�������9��h_�*��i�u�������L�ԓ�\9��C1��*��
�d�f�u�8�3���P���F��G1�*���f�d�%�u�j�u����&����|��[�����`�
�g�s�5�2�(���I����R��Q��@ۊ�g�u�u�:�;�%�2ߑ�����l ��\�����_�u�u�8��o����M¹��Z�_�����u�!�%�d��(�D���	���R��X ��*���
�|�0�&�w�m�L���YӒ��lW��Q��Eي�d�i�u����8���H�ӓ�l��^ �����l�
�d�g�w�}�W������]ǻN�����a�3�
�d��o�K�������@T��B1�F���u�'�;�!�?�o����IĹ��]ǻN�����b�1�8�'�6����K����Z���*���d�3�
�e�f�-�W���Y����Z9��h_�����e�b�%�|�]�}�W���&�ѓ�F9��1��U��}�8�
�d�1��D܁�J����lV�� 1�����d�
�f�n�w�}����H˹��lT��h�I���!�%�d�
�2��D������^��1����e�|�_�u�w�0�(�������9��R������-� �
�8�4����&����CW�N�����u�f�n�u�w�)��������9��R�����9�=�
�
�8�4����&����CW�N�Dʱ�"�!�u�|�]�}�W���&�֓�F9��1��U��3�
��-�"���������Q��G_��F���d�1�"�!�w�t�}���Y����W��B1�L���u�h�3�
��%����&����]��B1�@���}�e�1�"�#�}�D��Y����^��1��*��
�d�i�u���$����ԓ�\9��C1��*��
�d�g�u�w�}�������9F���*���3�
�g�
�e�a�Wǰ�����l ��_�����'�;�!�=�c�;�(��&���9F���*���3�
�a�
�e�a�Wǰ�����l ��]�����'�;�!�=�b�;�(��&���9F���*���1�8�'�4��(�F��&���F��Z��*���3�
�e�g�'�}��������ZR��1��*��m�%�|�_�w�}����L���� R��G\��H���8�
�f�3��o�(������^��1��*��
�g�n�u�w�)���&����W��N�U·�:�
��,�"��B߁�����l��N������e� �
�c����H����l�N����
� �m�b�'�}�J�������U��[��Gʺ�u�8�
�
�"�e�F���P���F��G1�*���m�d�%�u�j�W�W���Y�ƭ�l��D��Ҋ��"�0�u�#�-�D���&����CT�N��R��u�9�0�_�w�}�W���	����@��AV��N���u�!�%�g�1��Oہ�K�����E�����b�
�g�:�w�2��������9��UךU���8�
�e�3��o�(��E�ƪ�l��{:��:���d�d�<�
�/��(ށ�����l��N�Dʱ�"�!�u�|�]�}�W���&�ד�F9��1��U��_�u�u�u�w�0�(�������9�������8�
�m�3��m�(��I���W����ߊu�u�u�u�:��G���&����CW��N�����f�
� �c�f�-�W��Q����l��N!��*���
� �f�`�'�}�W�������)��h_�*���g�d�%�|�]�}�W���&�Փ�V��P�����d�`�%�u�j�u����&�ѓ�F9��]��Gʴ�1�!�%�<�>��A���&����l��d��Uʡ�%�f�
� �f�i�(��E����\��DX�� ��f�
�g�:�w�2����&����T��G\����u�8�
�m�1��F���	���N��C��M���
�e�c�%�w�/�����ޓ�F9��^��G��u�u�!�%�d�;�(��&���F�N�����&�2�0�}��%�"�������P��^ �����
�
� �b�n�-�^���
����WN��h�����#�a��|�w�1����[���F��G1�*���d�c�
�g�k�}�����ד�F9��Y��Gʺ�u�:�9�&��(�F��&���9F���*ߊ� �m�d�%�w�`�U���������Y�������g��#�l�F���&����e9��Q��Mӊ�g�u�u�<�9�9��������_��h_��U���0�w�w�_�w�}����@����l �� ]�����h�w�w�"�2�}����/����V��GZ��U���6�;�!�9�o��^ϻ�
���]ǻN�����
� �g�e�'�}�J�������A��\�U���u�8�
�
�2��E��B�����hV�� ��d�%�u�h�u�� ���Yے��lW��Q��Cۊ�a�h�4�
�8�.�(���&����_��^�����u�8�
�
�"�n�@���Y���D��_��]���
�d�3�
�a��C������]��[��C���9�0�w�w�]�}�W���&����^��N�U���4�%�4�d�#���������l��^�����:�g�|�_�w�}����&�ד�9��h_�B���u�h�w�w� �8�Wǲ�����l ��^�*��h�4�
�:�$�����I�Ʃ�@�L�U���!�%�<�<��(�F��&���F�N�����9�6��g�1��N؁�M����C9��Y������|�0�&�w�m�L���YӒ��l��1�*���d�b�
�g�k�}�G������_	��a1�����e�m�%�u�w�-�������� 9�������w�_�u�u�:��(�������T��N�U��u�=�;�}�8��(ہ�����9��S�����;�!�9�m��t����Y���9F���*���b�d�
� �f�n�(��E���F��R ������b�3�
�f�d����Y����\��h��F��u�9�0�w�u�W�W�������ZQ��B1�Fي�g�i�u�d�w�5��������9��h_�L���u�u�%�6�9�)����?����_��^�����u�8�
�
��n����Kƹ��Z�_�����u�9�6��f�;�(��&�����T�����g�
�|�0�$�}�G��Y����^��h�� ��l�%�u�h�u�� ���Yۊ��l0��B1�@���u�u�%�6�9�)����I�Ʃ�@�L�U���!�%�&�3��m�(��E���F��R �����d�
� �f�f�-�W���	����@��A]��\ʰ�&�u�e�n�2�9������